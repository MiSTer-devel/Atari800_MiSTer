
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(11 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 4095) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
        X"0b0b0b89",
        X"ad040b0b",
        X"0b0b0b0b",
        X"0b0b0b0b",
        X"0b0b0b0b",
        X"0b0b0b0b",
        X"0b0b0b0b",
        X"0b0b0b0b",
        X"0b0b0b0b",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"71fd0608",
        X"72830609",
        X"81058205",
        X"832b2a83",
        X"ffff0652",
        X"04000000",
        X"00000000",
        X"00000000",
        X"71fd0608",
        X"83ffff73",
        X"83060981",
        X"05820583",
        X"2b2b0906",
        X"7383ffff",
        X"0b0b0b0b",
        X"83a70400",
        X"72098105",
        X"72057373",
        X"09060906",
        X"73097306",
        X"070a8106",
        X"53510400",
        X"00000000",
        X"00000000",
        X"72722473",
        X"732e0753",
        X"51040000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"71737109",
        X"71068106",
        X"30720a10",
        X"0a720a10",
        X"0a31050a",
        X"81065151",
        X"53510400",
        X"00000000",
        X"72722673",
        X"732e0753",
        X"51040000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"0b0b0b88",
        X"bc040000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"720a722b",
        X"0a535104",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"72729f06",
        X"0981050b",
        X"0b0b889f",
        X"05040000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"72722aff",
        X"739f062a",
        X"0974090a",
        X"8106ff05",
        X"06075351",
        X"04000000",
        X"00000000",
        X"00000000",
        X"71715351",
        X"020d0406",
        X"73830609",
        X"81058205",
        X"832b0b2b",
        X"0772fc06",
        X"0c515104",
        X"00000000",
        X"72098105",
        X"72050970",
        X"81050906",
        X"0a810653",
        X"51040000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"72098105",
        X"72050970",
        X"81050906",
        X"0a098106",
        X"53510400",
        X"00000000",
        X"00000000",
        X"00000000",
        X"71098105",
        X"52040000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"72720981",
        X"05055351",
        X"04000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"72097206",
        X"73730906",
        X"07535104",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"71fc0608",
        X"72830609",
        X"81058305",
        X"1010102a",
        X"81ff0652",
        X"04000000",
        X"00000000",
        X"00000000",
        X"71fc0608",
        X"0b0b80e7",
        X"a4738306",
        X"10100508",
        X"060b0b0b",
        X"88a20400",
        X"00000000",
        X"00000000",
        X"0b0b0b88",
        X"ff040000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"0b0b0b88",
        X"d8040000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"72097081",
        X"0509060a",
        X"8106ff05",
        X"70547106",
        X"73097274",
        X"05ff0506",
        X"07515151",
        X"04000000",
        X"72097081",
        X"0509060a",
        X"098106ff",
        X"05705471",
        X"06730972",
        X"7405ff05",
        X"06075151",
        X"51040000",
        X"05ff0504",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"810b80ea",
        X"bc0c5104",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00007181",
        X"05520400",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000284",
        X"05721010",
        X"05520400",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00007171",
        X"05ff0571",
        X"5351020d",
        X"04000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"10101010",
        X"10101010",
        X"10101010",
        X"10101010",
        X"10101010",
        X"10101010",
        X"10101010",
        X"10101053",
        X"51047381",
        X"ff067383",
        X"06098105",
        X"83051010",
        X"102b0772",
        X"fc060c51",
        X"51043c04",
        X"72728072",
        X"8106ff05",
        X"09720605",
        X"71105272",
        X"0a100a53",
        X"72ed3851",
        X"51535104",
        X"83e08008",
        X"83e08408",
        X"83e08808",
        X"757580e5",
        X"c12d5050",
        X"83e08008",
        X"5683e088",
        X"0c83e084",
        X"0c83e080",
        X"0c510483",
        X"e0800883",
        X"e0840883",
        X"e0880875",
        X"7580e580",
        X"2d505083",
        X"e0800856",
        X"83e0880c",
        X"83e0840c",
        X"83e0800c",
        X"51040000",
        X"800489aa",
        X"0489aa0b",
        X"80decd04",
        X"fd3d0d75",
        X"705254af",
        X"b93f83e0",
        X"80081453",
        X"72742e92",
        X"38ff1370",
        X"33535371",
        X"af2e0981",
        X"06ee3881",
        X"13537283",
        X"e0800c85",
        X"3d0d04fd",
        X"3d0d7577",
        X"70535454",
        X"c73f83e0",
        X"8008732e",
        X"a13883e0",
        X"80087331",
        X"52ff1252",
        X"71ff2e8f",
        X"38727081",
        X"05543374",
        X"70810556",
        X"34eb39ff",
        X"14548074",
        X"34853d0d",
        X"04803d0d",
        X"7251ff90",
        X"3f823d0d",
        X"047183e0",
        X"800c0480",
        X"3d0d7251",
        X"80713481",
        X"0bbc120c",
        X"800b80c0",
        X"120c823d",
        X"0d04800b",
        X"83e2c008",
        X"248a38b6",
        X"8a3fff0b",
        X"83e2c00c",
        X"800b83e0",
        X"800c04ff",
        X"3d0d7352",
        X"83e09c08",
        X"722e8d38",
        X"d93f7151",
        X"96a03f71",
        X"83e09c0c",
        X"833d0d04",
        X"f43d0d7e",
        X"60625c5a",
        X"55805681",
        X"54bc1508",
        X"762e0981",
        X"06819138",
        X"7451c83f",
        X"7958757a",
        X"2580f738",
        X"83e2f008",
        X"70892a57",
        X"83ff0678",
        X"84807231",
        X"56565773",
        X"78258338",
        X"73557583",
        X"e2c0082e",
        X"8438ff82",
        X"3f83e2c0",
        X"088025a6",
        X"3875892b",
        X"5198dc3f",
        X"83e2f008",
        X"8f3dfc11",
        X"555c5481",
        X"52f81b51",
        X"96c63f76",
        X"1483e2f0",
        X"0c7583e2",
        X"c00c7453",
        X"76527851",
        X"b4b43f83",
        X"e0800883",
        X"e2f00816",
        X"83e2f00c",
        X"78763176",
        X"1b5b5956",
        X"778024ff",
        X"8b38617a",
        X"710c5475",
        X"5475802e",
        X"83388154",
        X"7383e080",
        X"0c8e3d0d",
        X"04fc3d0d",
        X"fe943f76",
        X"51fea83f",
        X"863dfc05",
        X"53785277",
        X"5195e93f",
        X"7975710c",
        X"5483e080",
        X"085483e0",
        X"8008802e",
        X"83388154",
        X"7383e080",
        X"0c863d0d",
        X"04fe3d0d",
        X"7583e2c0",
        X"08535380",
        X"72248938",
        X"71732e84",
        X"38fdcf3f",
        X"7451fde3",
        X"3f725197",
        X"ae3f83e0",
        X"80085283",
        X"e0800880",
        X"2e833881",
        X"527183e0",
        X"800c843d",
        X"0d04803d",
        X"0d7280c0",
        X"110883e0",
        X"800c5182",
        X"3d0d0480",
        X"3d0d72bc",
        X"110883e0",
        X"800c5182",
        X"3d0d0480",
        X"c40b83e0",
        X"800c04fd",
        X"3d0d7577",
        X"71547053",
        X"5553ab8a",
        X"3f82c813",
        X"08bc150c",
        X"82c01308",
        X"80c0150c",
        X"fce43f73",
        X"5193ab3f",
        X"7383e09c",
        X"0c83e080",
        X"085383e0",
        X"8008802e",
        X"83388153",
        X"7283e080",
        X"0c853d0d",
        X"04fd3d0d",
        X"75775553",
        X"fcb83f72",
        X"802ea538",
        X"bc130852",
        X"7351aa94",
        X"3f83e080",
        X"088f3877",
        X"527251ff",
        X"9a3f83e0",
        X"8008538a",
        X"3982cc13",
        X"0853d839",
        X"81537283",
        X"e0800c85",
        X"3d0d04fe",
        X"3d0dff0b",
        X"83e2c00c",
        X"7483e0a0",
        X"0c7583e2",
        X"bc0cb0e8",
        X"3f83e080",
        X"0881ff06",
        X"52815371",
        X"993883e2",
        X"d8518e94",
        X"3f83e080",
        X"085283e0",
        X"8008802e",
        X"83387252",
        X"71537283",
        X"e0800c84",
        X"3d0d04fa",
        X"3d0d787a",
        X"82c41208",
        X"82c41208",
        X"70722459",
        X"56565757",
        X"73732e09",
        X"81069138",
        X"80c01652",
        X"80c01751",
        X"a8853f83",
        X"e0800855",
        X"7483e080",
        X"0c883d0d",
        X"04f63d0d",
        X"7c5b807b",
        X"715c5457",
        X"7a772e8c",
        X"38811a82",
        X"cc140854",
        X"5a72f638",
        X"805980d9",
        X"397a5481",
        X"5780707b",
        X"7b315a57",
        X"55ff1853",
        X"74732580",
        X"c13882cc",
        X"14085273",
        X"51ff8c3f",
        X"800b83e0",
        X"800825a1",
        X"3882cc14",
        X"0882cc11",
        X"0882cc16",
        X"0c7482cc",
        X"120c5375",
        X"802e8638",
        X"7282cc17",
        X"0c725480",
        X"577382cc",
        X"15088117",
        X"575556ff",
        X"b8398119",
        X"59800bff",
        X"1b545478",
        X"73258338",
        X"81547681",
        X"32707506",
        X"515372ff",
        X"90388c3d",
        X"0d04f73d",
        X"0d7b7d5a",
        X"5a82d052",
        X"83e2bc08",
        X"5180d3fc",
        X"3f83e080",
        X"0857f9da",
        X"3f795283",
        X"e2c45195",
        X"b53f83e0",
        X"80085480",
        X"5383e080",
        X"08732e09",
        X"81068283",
        X"3883e0a0",
        X"080b0b80",
        X"e8dc5370",
        X"5256a7c2",
        X"3f0b0b80",
        X"e8dc5280",
        X"c01651a7",
        X"b53f75bc",
        X"170c7382",
        X"c0170c81",
        X"0b82c417",
        X"0c810b82",
        X"c8170c73",
        X"82cc170c",
        X"ff1782d0",
        X"17555781",
        X"913983e0",
        X"ac337082",
        X"2a708106",
        X"51545572",
        X"81803874",
        X"812a8106",
        X"587780f6",
        X"3874842a",
        X"810682c4",
        X"150c83e0",
        X"ac338106",
        X"82c8150c",
        X"79527351",
        X"a6dc3f73",
        X"51a6f33f",
        X"83e08008",
        X"1453af73",
        X"70810555",
        X"3472bc15",
        X"0c83e0ad",
        X"527251a6",
        X"bd3f83e0",
        X"a40882c0",
        X"150c83e0",
        X"ba5280c0",
        X"1451a6aa",
        X"3f78802e",
        X"8d387351",
        X"782d83e0",
        X"8008802e",
        X"99387782",
        X"cc150c75",
        X"802e8638",
        X"7382cc17",
        X"0c7382d0",
        X"15ff1959",
        X"55567680",
        X"2e9b3883",
        X"e0a45283",
        X"e2c45194",
        X"ab3f83e0",
        X"80088a38",
        X"83e0ad33",
        X"5372fed2",
        X"3878802e",
        X"893883e0",
        X"a00851fc",
        X"b83f83e0",
        X"a0085372",
        X"83e0800c",
        X"8b3d0d04",
        X"ff3d0d80",
        X"527351fd",
        X"b53f833d",
        X"0d04f03d",
        X"0d627052",
        X"54f6893f",
        X"83e08008",
        X"7453873d",
        X"70535555",
        X"f6a93ff7",
        X"893f7351",
        X"d33f6353",
        X"745283e0",
        X"800851fa",
        X"b83f923d",
        X"0d047183",
        X"e0800c04",
        X"80c01283",
        X"e0800c04",
        X"803d0d72",
        X"82c01108",
        X"83e0800c",
        X"51823d0d",
        X"04803d0d",
        X"7282cc11",
        X"0883e080",
        X"0c51823d",
        X"0d04803d",
        X"0d7282c4",
        X"110883e0",
        X"800c5182",
        X"3d0d04f9",
        X"3d0d7983",
        X"e0900857",
        X"57817727",
        X"81963876",
        X"88170827",
        X"818e3875",
        X"33557482",
        X"2e893874",
        X"832eb338",
        X"80fe3974",
        X"54761083",
        X"fe065376",
        X"882a8c17",
        X"08055289",
        X"3dfc0551",
        X"ab963f83",
        X"e0800880",
        X"df38029d",
        X"0533893d",
        X"3371882b",
        X"07565680",
        X"d1398454",
        X"76822b83",
        X"fc065376",
        X"872a8c17",
        X"08055289",
        X"3dfc0551",
        X"aae63f83",
        X"e08008b0",
        X"38029f05",
        X"33028405",
        X"9e053371",
        X"982b7190",
        X"2b07028c",
        X"059d0533",
        X"70882b72",
        X"078d3d33",
        X"7180ffff",
        X"fe800607",
        X"51525357",
        X"58568339",
        X"81557483",
        X"e0800c89",
        X"3d0d04fb",
        X"3d0d83e0",
        X"9008fe19",
        X"881208fe",
        X"05555654",
        X"80567473",
        X"278d3882",
        X"14337571",
        X"29941608",
        X"05575375",
        X"83e0800c",
        X"873d0d04",
        X"fc3d0d76",
        X"52800b83",
        X"e0900870",
        X"33515253",
        X"70832e09",
        X"81069138",
        X"95123394",
        X"13337198",
        X"2b71902b",
        X"07555551",
        X"9b12339a",
        X"13337188",
        X"2b077407",
        X"83e0800c",
        X"55863d0d",
        X"04fc3d0d",
        X"7683e090",
        X"08555580",
        X"75238815",
        X"08537281",
        X"2e883888",
        X"14087326",
        X"85388152",
        X"b2397290",
        X"38733352",
        X"71832e09",
        X"81068538",
        X"90140853",
        X"728c160c",
        X"72802e8d",
        X"387251fe",
        X"d63f83e0",
        X"80085285",
        X"39901408",
        X"52719016",
        X"0c805271",
        X"83e0800c",
        X"863d0d04",
        X"fa3d0d78",
        X"83e09008",
        X"71228105",
        X"7083ffff",
        X"06575457",
        X"5573802e",
        X"88389015",
        X"08537286",
        X"38835280",
        X"e739738f",
        X"06527180",
        X"da388113",
        X"90160c8c",
        X"15085372",
        X"9038830b",
        X"84172257",
        X"52737627",
        X"80c638bf",
        X"39821633",
        X"ff057484",
        X"2a065271",
        X"b2387251",
        X"fcb13f81",
        X"527183e0",
        X"800827a8",
        X"38835283",
        X"e0800888",
        X"1708279c",
        X"3883e080",
        X"088c160c",
        X"83e08008",
        X"51fdbc3f",
        X"83e08008",
        X"90160c73",
        X"75238052",
        X"7183e080",
        X"0c883d0d",
        X"04f23d0d",
        X"60626458",
        X"5e5b7533",
        X"5574a02e",
        X"09810688",
        X"38811670",
        X"4456ef39",
        X"62703356",
        X"5674af2e",
        X"09810684",
        X"38811643",
        X"800b881c",
        X"0c627033",
        X"5155749f",
        X"2691387a",
        X"51fdd23f",
        X"83e08008",
        X"56807d34",
        X"83813993",
        X"3d841c08",
        X"7058595f",
        X"8a55a076",
        X"70810558",
        X"34ff1555",
        X"74ff2e09",
        X"8106ef38",
        X"80705a5c",
        X"887f085f",
        X"5a7b811d",
        X"7081ff06",
        X"60137033",
        X"70af3270",
        X"30a07327",
        X"71802507",
        X"5151525b",
        X"535e5755",
        X"7480e738",
        X"76ae2e09",
        X"81068338",
        X"8155787a",
        X"27750755",
        X"74802e9f",
        X"38798832",
        X"703078ae",
        X"32703070",
        X"73079f2a",
        X"53515751",
        X"5675bb38",
        X"88598b5a",
        X"ffab3976",
        X"982b5574",
        X"80258738",
        X"80e6b417",
        X"3357ff9f",
        X"17557499",
        X"268938e0",
        X"177081ff",
        X"06585578",
        X"811a7081",
        X"ff067a13",
        X"535b5755",
        X"767534fe",
        X"f8397b1e",
        X"7f0c8055",
        X"76a02683",
        X"38815574",
        X"8b19347a",
        X"51fc823f",
        X"83e08008",
        X"80f538a0",
        X"547a2270",
        X"852b83e0",
        X"06545590",
        X"1b08527c",
        X"51a5a13f",
        X"83e08008",
        X"5783e080",
        X"08818138",
        X"7c335574",
        X"802e80f4",
        X"388b1d33",
        X"70832a70",
        X"81065156",
        X"5674b438",
        X"8b7d841d",
        X"0883e080",
        X"08595b5b",
        X"58ff1858",
        X"77ff2e9a",
        X"38797081",
        X"055b3379",
        X"7081055b",
        X"33717131",
        X"52565675",
        X"802ee238",
        X"86397580",
        X"2e96387a",
        X"51fbe53f",
        X"ff863983",
        X"e0800856",
        X"83e08008",
        X"b6388339",
        X"7656841b",
        X"088b1133",
        X"515574a7",
        X"388b1d33",
        X"70842a70",
        X"81065156",
        X"56748938",
        X"83569439",
        X"81569039",
        X"7c51fa94",
        X"3f83e080",
        X"08881c0c",
        X"fd813975",
        X"83e0800c",
        X"903d0d04",
        X"f83d0d7a",
        X"7c595782",
        X"5483fe53",
        X"77527651",
        X"a3e63f83",
        X"5683e080",
        X"0880ec38",
        X"81173377",
        X"3371882b",
        X"07565682",
        X"567482d4",
        X"d52e0981",
        X"0680d438",
        X"7554b653",
        X"77527651",
        X"a3ba3f83",
        X"e0800898",
        X"38811733",
        X"77337188",
        X"2b0783e0",
        X"80085256",
        X"56748182",
        X"c62eac38",
        X"825480d2",
        X"53775276",
        X"51a3913f",
        X"83e08008",
        X"98388117",
        X"33773371",
        X"882b0783",
        X"e0800852",
        X"56567481",
        X"82c62e83",
        X"38815675",
        X"83e0800c",
        X"8a3d0d04",
        X"eb3d0d67",
        X"5a800b83",
        X"e0900ca2",
        X"b33f83e0",
        X"80088106",
        X"55825674",
        X"83ef3874",
        X"75538f3d",
        X"70535759",
        X"feca3f83",
        X"e0800881",
        X"ff065776",
        X"812e0981",
        X"0680d438",
        X"905483be",
        X"53745275",
        X"51a2a53f",
        X"83e08008",
        X"80c9388f",
        X"3d335574",
        X"802e80c9",
        X"3802bf05",
        X"33028405",
        X"be053371",
        X"982b7190",
        X"2b07028c",
        X"05bd0533",
        X"70882b72",
        X"07953d33",
        X"71077058",
        X"7b575e52",
        X"5e575957",
        X"fdee3f83",
        X"e0800881",
        X"ff065776",
        X"832e0981",
        X"06863881",
        X"5682f239",
        X"76802e86",
        X"38865682",
        X"e839a454",
        X"8d537852",
        X"7551a1bc",
        X"3f815683",
        X"e0800882",
        X"d43802be",
        X"05330284",
        X"05bd0533",
        X"71882b07",
        X"595d77ab",
        X"380280ce",
        X"05330284",
        X"0580cd05",
        X"3371982b",
        X"71902b07",
        X"973d3370",
        X"882b7207",
        X"02940580",
        X"cb053371",
        X"0754525e",
        X"57595602",
        X"b7053378",
        X"71290288",
        X"05b60533",
        X"028c05b5",
        X"05337188",
        X"2b07701d",
        X"707f8c05",
        X"0c5f5957",
        X"595d8e3d",
        X"33821b34",
        X"02b90533",
        X"903d3371",
        X"882b075a",
        X"5c78841b",
        X"2302bb05",
        X"33028405",
        X"ba053371",
        X"882b0756",
        X"5c74ab38",
        X"0280ca05",
        X"33028405",
        X"80c90533",
        X"71982b71",
        X"902b0796",
        X"3d337088",
        X"2b720702",
        X"940580c7",
        X"05337107",
        X"51525357",
        X"5e5c7476",
        X"31783179",
        X"842a903d",
        X"33547171",
        X"31535656",
        X"80c4e13f",
        X"83e08008",
        X"82057088",
        X"1c0c83e0",
        X"8008e08a",
        X"05565674",
        X"83dffe26",
        X"83388257",
        X"83fff676",
        X"27853883",
        X"57893986",
        X"5676802e",
        X"80db3876",
        X"7a347683",
        X"2e098106",
        X"b0380280",
        X"d6053302",
        X"840580d5",
        X"05337198",
        X"2b71902b",
        X"07993d33",
        X"70882b72",
        X"07029405",
        X"80d30533",
        X"71077f90",
        X"050c525e",
        X"57585686",
        X"39771b90",
        X"1b0c841a",
        X"228c1b08",
        X"1971842a",
        X"05941c0c",
        X"5d800b81",
        X"1b347983",
        X"e0900c80",
        X"567583e0",
        X"800c973d",
        X"0d04e93d",
        X"0d83e090",
        X"08568554",
        X"75802e81",
        X"8238800b",
        X"81173499",
        X"3de01146",
        X"6a548a3d",
        X"705458ec",
        X"0551f6e5",
        X"3f83e080",
        X"085483e0",
        X"800880df",
        X"38893d33",
        X"5473802e",
        X"913802ab",
        X"05337084",
        X"2a810651",
        X"5574802e",
        X"86388354",
        X"80c13976",
        X"51f4893f",
        X"83e08008",
        X"a0170c02",
        X"bf053302",
        X"8405be05",
        X"3371982b",
        X"71902b07",
        X"028c05bd",
        X"05337088",
        X"2b720795",
        X"3d337107",
        X"9c1c0c52",
        X"78981b0c",
        X"53565957",
        X"810b8117",
        X"34745473",
        X"83e0800c",
        X"993d0d04",
        X"f53d0d7d",
        X"7f617283",
        X"e090085a",
        X"5d5d595c",
        X"807b0c85",
        X"5775802e",
        X"81e03881",
        X"16338106",
        X"55845774",
        X"802e81d2",
        X"38913974",
        X"81173486",
        X"39800b81",
        X"17348157",
        X"81c0399c",
        X"16089817",
        X"08315574",
        X"78278338",
        X"74587780",
        X"2e81a938",
        X"98160870",
        X"83ff0656",
        X"577480cf",
        X"38821633",
        X"ff057789",
        X"2a067081",
        X"ff065a55",
        X"78a03876",
        X"8738a016",
        X"08558d39",
        X"a4160851",
        X"f0e93f83",
        X"e0800855",
        X"817527ff",
        X"a83874a4",
        X"170ca416",
        X"0851f283",
        X"3f83e080",
        X"085583e0",
        X"8008802e",
        X"ff893883",
        X"e0800819",
        X"a8170c98",
        X"160883ff",
        X"06848071",
        X"31515577",
        X"75278338",
        X"77557483",
        X"ffff0654",
        X"98160883",
        X"ff0653a8",
        X"16085279",
        X"577b8338",
        X"7b577651",
        X"9be23f83",
        X"e08008fe",
        X"d0389816",
        X"08159817",
        X"0c741a78",
        X"76317c08",
        X"177d0c59",
        X"5afed339",
        X"80577683",
        X"e0800c8d",
        X"3d0d04fa",
        X"3d0d7883",
        X"e0900855",
        X"56855573",
        X"802e81e1",
        X"38811433",
        X"81065384",
        X"5572802e",
        X"81d3389c",
        X"14085372",
        X"76278338",
        X"72569814",
        X"0857800b",
        X"98150c75",
        X"802e81b7",
        X"38821433",
        X"70892b56",
        X"5376802e",
        X"b5387452",
        X"ff1651bf",
        X"e33f83e0",
        X"8008ff18",
        X"76547053",
        X"5853bfd4",
        X"3f83e080",
        X"08732696",
        X"38743070",
        X"78067098",
        X"170c7771",
        X"31a41708",
        X"52585153",
        X"8939a014",
        X"0870a416",
        X"0c537476",
        X"27b93872",
        X"51eed83f",
        X"83e08008",
        X"53810b83",
        X"e0800827",
        X"8b388814",
        X"0883e080",
        X"08268838",
        X"800b8115",
        X"34b03983",
        X"e08008a4",
        X"150c9814",
        X"08159815",
        X"0c757531",
        X"56c43998",
        X"14081670",
        X"98160c73",
        X"5256efc7",
        X"3f83e080",
        X"088c3883",
        X"e0800881",
        X"15348155",
        X"94398214",
        X"33ff0576",
        X"892a0683",
        X"e0800805",
        X"a8150c80",
        X"557483e0",
        X"800c883d",
        X"0d04ef3d",
        X"0d635685",
        X"5583e090",
        X"08802e80",
        X"d238933d",
        X"f4058417",
        X"0c645388",
        X"3d705376",
        X"5257f1d1",
        X"3f83e080",
        X"085583e0",
        X"8008b438",
        X"883d3354",
        X"73802ea1",
        X"3802a705",
        X"3370842a",
        X"70810651",
        X"55558355",
        X"73802e97",
        X"387651ee",
        X"f73f83e0",
        X"80088817",
        X"0c7551ef",
        X"a83f83e0",
        X"80085574",
        X"83e0800c",
        X"933d0d04",
        X"e43d0d6e",
        X"a13d0840",
        X"5e855683",
        X"e0900880",
        X"2e848538",
        X"9e3df405",
        X"841f0c7e",
        X"98387d51",
        X"eef73f83",
        X"e0800856",
        X"83ee3981",
        X"4181f639",
        X"834181f1",
        X"39933d7f",
        X"96054159",
        X"807f8295",
        X"055e5675",
        X"6081ff05",
        X"34834190",
        X"1e08762e",
        X"81d338a0",
        X"547d2270",
        X"852b83e0",
        X"06545890",
        X"1e085278",
        X"5197ed3f",
        X"83e08008",
        X"4183e080",
        X"08ffb838",
        X"78335c7b",
        X"802effb4",
        X"388b1933",
        X"70bf0671",
        X"81065243",
        X"5574802e",
        X"80de387b",
        X"81bf0655",
        X"748f2480",
        X"d3389a19",
        X"33557480",
        X"cb38f31d",
        X"70585d81",
        X"56758b2e",
        X"09810685",
        X"388e568b",
        X"39759a2e",
        X"09810683",
        X"389c5678",
        X"16707081",
        X"05523371",
        X"33811a82",
        X"1a5f5b52",
        X"5b557486",
        X"38797734",
        X"853980df",
        X"7734777b",
        X"57577aa0",
        X"2e098106",
        X"c0388156",
        X"7b81e532",
        X"7030709f",
        X"2a515155",
        X"7bae2e93",
        X"3874802e",
        X"8e386183",
        X"2a708106",
        X"51557480",
        X"2e97387d",
        X"51ede13f",
        X"83e08008",
        X"4183e080",
        X"08873890",
        X"1e08feaf",
        X"38806034",
        X"75802e88",
        X"387c527f",
        X"518f933f",
        X"60802e86",
        X"38800b90",
        X"1f0c6056",
        X"60832e85",
        X"386081d0",
        X"38891f57",
        X"901e0880",
        X"2e81a838",
        X"80567816",
        X"70335155",
        X"74a02ea0",
        X"3874852e",
        X"09810684",
        X"3881e555",
        X"74777081",
        X"05593481",
        X"167081ff",
        X"06575587",
        X"7627d738",
        X"88193355",
        X"74a02ea9",
        X"38ae7770",
        X"81055934",
        X"88567816",
        X"70335155",
        X"74a02e95",
        X"38747770",
        X"81055934",
        X"81167081",
        X"ff065755",
        X"8a7627e2",
        X"388b1933",
        X"7f880534",
        X"9f19339e",
        X"1a337198",
        X"2b71902b",
        X"079d1c33",
        X"70882b72",
        X"079c1e33",
        X"7107640c",
        X"52991d33",
        X"981e3371",
        X"882b0753",
        X"51535759",
        X"56747f84",
        X"05239719",
        X"33961a33",
        X"71882b07",
        X"5656747f",
        X"86052380",
        X"77347d51",
        X"ebf23f83",
        X"e0800883",
        X"32703070",
        X"72079f2c",
        X"83e08008",
        X"06525656",
        X"961f3355",
        X"748a3889",
        X"1f52961f",
        X"518d9f3f",
        X"7583e080",
        X"0c9e3d0d",
        X"04f43d0d",
        X"7e8f3dec",
        X"11565658",
        X"9053f015",
        X"527751e0",
        X"d43f83e0",
        X"800880d6",
        X"3878902e",
        X"09810680",
        X"cd3802ab",
        X"053380ea",
        X"c40b80ea",
        X"c4335758",
        X"568c3974",
        X"762e8a38",
        X"84177033",
        X"565774f3",
        X"38763370",
        X"57557480",
        X"2eac3882",
        X"1722708a",
        X"2b903dec",
        X"05567055",
        X"56569680",
        X"0a527751",
        X"e0833f83",
        X"e0800886",
        X"3878752e",
        X"85388056",
        X"85398117",
        X"33567583",
        X"e0800c8e",
        X"3d0d04fc",
        X"3d0d7670",
        X"52558ca6",
        X"3f83e080",
        X"0815ff05",
        X"5473752e",
        X"8e387333",
        X"5372ae2e",
        X"8638ff14",
        X"54ef3977",
        X"52811451",
        X"8bbe3f83",
        X"e0800830",
        X"7083e080",
        X"08078025",
        X"83e0800c",
        X"53863d0d",
        X"04fc3d0d",
        X"76705255",
        X"e6f03f83",
        X"e0800854",
        X"815383e0",
        X"800880c1",
        X"387451e6",
        X"b33f83e0",
        X"800880e8",
        X"e05383e0",
        X"80085253",
        X"ff913f83",
        X"e08008a1",
        X"3880e8e4",
        X"527251ff",
        X"823f83e0",
        X"80089238",
        X"80e8e852",
        X"7251fef3",
        X"3f83e080",
        X"08802e83",
        X"38815473",
        X"537283e0",
        X"800c863d",
        X"0d04fc3d",
        X"0d767052",
        X"55e68f3f",
        X"83e08008",
        X"54815383",
        X"e0800880",
        X"d1387451",
        X"e5d23f83",
        X"e0800880",
        X"e8e05383",
        X"e0800852",
        X"53feb03f",
        X"83e08008",
        X"b13880e8",
        X"e4527251",
        X"fea13f83",
        X"e08008a2",
        X"3880e8e8",
        X"527251fe",
        X"923f83e0",
        X"80089338",
        X"83e39808",
        X"527251fe",
        X"823f83e0",
        X"8008802e",
        X"83388154",
        X"73537283",
        X"e0800c86",
        X"3d0d04fd",
        X"3d0d7570",
        X"5254e59e",
        X"3f815383",
        X"e0800898",
        X"387351e4",
        X"e73f83e3",
        X"88085283",
        X"e0800851",
        X"fdc93f83",
        X"e0800853",
        X"7283e080",
        X"0c853d0d",
        X"04df3d0d",
        X"a43d0870",
        X"525edb85",
        X"3f83e080",
        X"0833953d",
        X"56547396",
        X"3880ebcc",
        X"52745189",
        X"ad3f9a39",
        X"7d527851",
        X"de8d3f84",
        X"ca397d51",
        X"daeb3f83",
        X"e0800852",
        X"7451da9b",
        X"3f804380",
        X"42804180",
        X"4083e390",
        X"0852943d",
        X"70525de0",
        X"f53f83e0",
        X"80085980",
        X"0b83e080",
        X"08555b83",
        X"e080087b",
        X"2e943881",
        X"1b74525b",
        X"e3f73f83",
        X"e0800854",
        X"83e08008",
        X"ee38805a",
        X"ff5f7909",
        X"709f2c7b",
        X"065b547a",
        X"7a248438",
        X"ff1b5af6",
        X"1a700970",
        X"9f2c7206",
        X"7bff125a",
        X"5a525555",
        X"80752595",
        X"387651e3",
        X"bc3f83e0",
        X"800876ff",
        X"18585557",
        X"738024ed",
        X"38747f2e",
        X"8638a19b",
        X"3f745f78",
        X"ff1b7058",
        X"5d58807a",
        X"25953877",
        X"51e3923f",
        X"83e08008",
        X"76ff1858",
        X"55587380",
        X"24ed3880",
        X"0b83e7c0",
        X"0c800b83",
        X"e7ec0c80",
        X"e8ec518d",
        X"ac3f8180",
        X"0b83e7ec",
        X"0c80e8f4",
        X"518d9e3f",
        X"a80b83e7",
        X"c00c7680",
        X"2e80e438",
        X"83e7c008",
        X"77793270",
        X"30707207",
        X"80257087",
        X"2b83e7ec",
        X"0c515678",
        X"535656e2",
        X"c93f83e0",
        X"8008802e",
        X"883880e8",
        X"fc518ce5",
        X"3f7651e2",
        X"8b3f83e0",
        X"80085280",
        X"ea8c518c",
        X"d43f7651",
        X"e2933f83",
        X"e0800883",
        X"e7c00855",
        X"57757425",
        X"8638a816",
        X"56f73975",
        X"83e7c00c",
        X"86f07624",
        X"ff983887",
        X"980b83e7",
        X"c00c7780",
        X"2eb13877",
        X"51e1c93f",
        X"83e08008",
        X"785255e1",
        X"e93f80e9",
        X"845483e0",
        X"80088d38",
        X"87398076",
        X"3481ea39",
        X"80e8b454",
        X"74537352",
        X"80e98851",
        X"8bf33f80",
        X"5480e990",
        X"518bea3f",
        X"81145473",
        X"a82e0981",
        X"06ef3886",
        X"8da0519d",
        X"8f3f8052",
        X"903d7052",
        X"58b18f3f",
        X"83527751",
        X"b1883f62",
        X"81ab3861",
        X"802e8197",
        X"387b5473",
        X"ff2e9638",
        X"78802e81",
        X"86387851",
        X"e0ef3f83",
        X"e08008ff",
        X"155559e7",
        X"3978802e",
        X"80f13878",
        X"51e0eb3f",
        X"83e08008",
        X"802efc90",
        X"387851e0",
        X"b33f83e0",
        X"80085280",
        X"e8dc5184",
        X"823f83e0",
        X"8008bb38",
        X"7c5185ba",
        X"3f83e080",
        X"08ff0555",
        X"800b83e0",
        X"80082580",
        X"c838a33d",
        X"7505c405",
        X"70585676",
        X"33ff1858",
        X"5473af2e",
        X"fec43874",
        X"ff16ff18",
        X"58565473",
        X"8024e838",
        X"a4397851",
        X"dfdc3f83",
        X"e0800852",
        X"7c5184da",
        X"3f933981",
        X"549e397f",
        X"10608829",
        X"057a0561",
        X"055afbf6",
        X"3962802e",
        X"fbb73880",
        X"527751af",
        X"cd3f8054",
        X"7383e080",
        X"0ca33d0d",
        X"04803d0d",
        X"9088b833",
        X"7081ff06",
        X"70842a81",
        X"32708106",
        X"51515151",
        X"70802e8d",
        X"38a80b90",
        X"88b834b8",
        X"0b9088b8",
        X"347083e0",
        X"800c823d",
        X"0d04803d",
        X"0d9088b8",
        X"337081ff",
        X"0670852a",
        X"81327081",
        X"06515151",
        X"5170802e",
        X"8d38980b",
        X"9088b834",
        X"b80b9088",
        X"b8347083",
        X"e0800c82",
        X"3d0d0493",
        X"0b9088bc",
        X"34ff0b90",
        X"88a83404",
        X"ff3d0d02",
        X"8f053352",
        X"800b9088",
        X"bc348a51",
        X"9ab63fdf",
        X"3f80f80b",
        X"9088a034",
        X"800b9088",
        X"8834fa12",
        X"52719088",
        X"8034800b",
        X"90889834",
        X"71908890",
        X"349088b8",
        X"52807234",
        X"b8723483",
        X"3d0d0480",
        X"3d0d028b",
        X"05335170",
        X"9088b434",
        X"febf3f83",
        X"e0800880",
        X"2ef63882",
        X"3d0d0480",
        X"3d0d8439",
        X"a6c13ffe",
        X"d93f83e0",
        X"8008802e",
        X"f3389088",
        X"b4337081",
        X"ff0683e0",
        X"800c5182",
        X"3d0d0480",
        X"3d0da30b",
        X"9088bc34",
        X"ff0b9088",
        X"a8349088",
        X"b851a871",
        X"34b87134",
        X"823d0d04",
        X"803d0d90",
        X"88bc3370",
        X"982b7080",
        X"2583e080",
        X"0c515182",
        X"3d0d0480",
        X"3d0d9088",
        X"b8337081",
        X"ff067083",
        X"2a813270",
        X"81065151",
        X"51517080",
        X"2ee838b0",
        X"0b9088b8",
        X"34b80b90",
        X"88b83482",
        X"3d0d0480",
        X"3d0d9080",
        X"ac088106",
        X"83e0800c",
        X"823d0d04",
        X"fd3d0d75",
        X"77545480",
        X"73259438",
        X"73708105",
        X"55335280",
        X"e9945187",
        X"843fff13",
        X"53e93985",
        X"3d0d04fd",
        X"3d0d7577",
        X"53547333",
        X"51708938",
        X"71335170",
        X"802ea138",
        X"73337233",
        X"52537271",
        X"278538ff",
        X"51943970",
        X"73278538",
        X"81518b39",
        X"81148113",
        X"5354d339",
        X"80517083",
        X"e0800c85",
        X"3d0d04fd",
        X"3d0d7577",
        X"54547233",
        X"7081ff06",
        X"52527080",
        X"2ea33871",
        X"81ff0681",
        X"14ffbf12",
        X"53545270",
        X"99268938",
        X"a0127081",
        X"ff065351",
        X"71747081",
        X"055634d2",
        X"39807434",
        X"853d0d04",
        X"ffbd3d0d",
        X"80c63d08",
        X"52a53d70",
        X"5254ffb3",
        X"3f80c73d",
        X"0852853d",
        X"705253ff",
        X"a63f7252",
        X"7351fedf",
        X"3f80c53d",
        X"0d04fe3d",
        X"0d747653",
        X"53717081",
        X"05533351",
        X"70737081",
        X"05553470",
        X"f038843d",
        X"0d04fe3d",
        X"0d745280",
        X"72335253",
        X"70732e8d",
        X"38811281",
        X"14713353",
        X"545270f5",
        X"387283e0",
        X"800c843d",
        X"0d04f63d",
        X"0d7c7e60",
        X"625a5d5b",
        X"56805981",
        X"55853974",
        X"7a295574",
        X"527551ab",
        X"ab3f83e0",
        X"80087a27",
        X"ee387480",
        X"2e80dd38",
        X"74527551",
        X"ab963f83",
        X"e0800875",
        X"53765254",
        X"ab9a3f83",
        X"e080087a",
        X"53755256",
        X"aafe3f83",
        X"e0800879",
        X"30707b07",
        X"9f2a7077",
        X"80240751",
        X"51545572",
        X"873883e0",
        X"8008c538",
        X"768118b0",
        X"16555858",
        X"8974258b",
        X"38b71453",
        X"7a853880",
        X"d7145372",
        X"78348119",
        X"59ff9f39",
        X"8077348c",
        X"3d0d04f7",
        X"3d0d7b7d",
        X"7f620290",
        X"05bb0533",
        X"5759565a",
        X"5ab05872",
        X"8338a058",
        X"75707081",
        X"05523371",
        X"59545590",
        X"39807425",
        X"8e38ff14",
        X"77708105",
        X"59335454",
        X"72ef3873",
        X"ff155553",
        X"80732589",
        X"38775279",
        X"51782def",
        X"39753375",
        X"57537280",
        X"2e903872",
        X"52795178",
        X"2d757081",
        X"05573353",
        X"ed398b3d",
        X"0d04ee3d",
        X"0d646669",
        X"69707081",
        X"0552335b",
        X"4a5c5e5e",
        X"76802e82",
        X"f93876a5",
        X"2e098106",
        X"82e03880",
        X"70416770",
        X"70810552",
        X"33714a59",
        X"575f76b0",
        X"2e098106",
        X"8c387570",
        X"81055733",
        X"76485781",
        X"5fd01756",
        X"75892680",
        X"da387667",
        X"5c59805c",
        X"9339778a",
        X"2480c338",
        X"7b8a2918",
        X"7b708105",
        X"5d335a5c",
        X"d0197081",
        X"ff065858",
        X"897727a4",
        X"38ff9f19",
        X"7081ff06",
        X"ffa91b5a",
        X"51568576",
        X"279238ff",
        X"bf197081",
        X"ff065156",
        X"7585268a",
        X"38c91958",
        X"778025ff",
        X"b9387a47",
        X"7b407881",
        X"ff065776",
        X"80e42e80",
        X"e5387680",
        X"e424a738",
        X"7680d82e",
        X"81863876",
        X"80d82490",
        X"3876802e",
        X"81cc3876",
        X"a52e81b6",
        X"3881b939",
        X"7680e32e",
        X"818c3881",
        X"af397680",
        X"f52e9b38",
        X"7680f524",
        X"8b387680",
        X"f32e8181",
        X"38819939",
        X"7680f82e",
        X"80ca3881",
        X"8f39913d",
        X"70555780",
        X"538a5279",
        X"841b7108",
        X"535b56fc",
        X"813f7655",
        X"ab397984",
        X"1b710894",
        X"3d705b5b",
        X"525b5675",
        X"80258c38",
        X"753056ad",
        X"78340280",
        X"c1055776",
        X"5480538a",
        X"527551fb",
        X"d53f7755",
        X"7e54b839",
        X"913d7055",
        X"7780d832",
        X"70307080",
        X"25565158",
        X"56905279",
        X"841b7108",
        X"535b57fb",
        X"b13f7555",
        X"db397984",
        X"1b831233",
        X"545b5698",
        X"3979841b",
        X"7108575b",
        X"5680547f",
        X"537c527d",
        X"51fc9c3f",
        X"87397652",
        X"7d517c2d",
        X"66703358",
        X"810547fd",
        X"8339943d",
        X"0d047283",
        X"e0940c71",
        X"83e0980c",
        X"04fb3d0d",
        X"883d7070",
        X"84055208",
        X"57547553",
        X"83e09408",
        X"5283e098",
        X"0851fcc6",
        X"3f873d0d",
        X"04ff3d0d",
        X"73700853",
        X"51029305",
        X"33723470",
        X"08810571",
        X"0c833d0d",
        X"04fc3d0d",
        X"873d8811",
        X"557854be",
        X"cd5351fc",
        X"993f8052",
        X"873d51d1",
        X"3f863d0d",
        X"04fc3d0d",
        X"76557483",
        X"e39c082e",
        X"af388053",
        X"745187c6",
        X"3f83e080",
        X"0881ff06",
        X"ff147081",
        X"ff067230",
        X"709f2a51",
        X"52555354",
        X"72802e84",
        X"3871dd38",
        X"73fe3874",
        X"83e39c0c",
        X"863d0d04",
        X"ff3d0dff",
        X"0b83e39c",
        X"0c84a53f",
        X"8151878a",
        X"3f83e080",
        X"0881ff06",
        X"5271ee38",
        X"81d33f71",
        X"83e0800c",
        X"833d0d04",
        X"fc3d0d76",
        X"028405a2",
        X"05220288",
        X"05a60522",
        X"7a545555",
        X"55ff823f",
        X"72802ea0",
        X"3883e3b0",
        X"14337570",
        X"81055734",
        X"81147083",
        X"ffff06ff",
        X"157083ff",
        X"ff065652",
        X"5552dd39",
        X"800b83e0",
        X"800c863d",
        X"0d04fc3d",
        X"0d76787a",
        X"11565355",
        X"80537174",
        X"2e933874",
        X"13517033",
        X"83e3b013",
        X"34811281",
        X"145452ea",
        X"39800b83",
        X"e0800c86",
        X"3d0d04fd",
        X"3d0d9054",
        X"83e39c08",
        X"5186f93f",
        X"83e08008",
        X"81ff06ff",
        X"15713071",
        X"30707307",
        X"9f2a729f",
        X"2a065255",
        X"52555372",
        X"db38853d",
        X"0d04803d",
        X"0d83e3a8",
        X"081083e3",
        X"a0080790",
        X"80a80c82",
        X"3d0d0480",
        X"0b83e3a8",
        X"0ce43f04",
        X"810b83e3",
        X"a80cdb3f",
        X"04ed3f04",
        X"7183e3a4",
        X"0c04803d",
        X"0d8051f4",
        X"3f810b83",
        X"e3a80c81",
        X"0b83e3a0",
        X"0cffbb3f",
        X"823d0d04",
        X"803d0d72",
        X"30707407",
        X"802583e3",
        X"a00c51ff",
        X"a53f823d",
        X"0d04803d",
        X"0d028b05",
        X"339080a4",
        X"0c9080a8",
        X"08708106",
        X"515170f5",
        X"389080a4",
        X"087081ff",
        X"0683e080",
        X"0c51823d",
        X"0d04803d",
        X"0d81ff51",
        X"d13f83e0",
        X"800881ff",
        X"0683e080",
        X"0c823d0d",
        X"04803d0d",
        X"73902b73",
        X"079080b4",
        X"0c823d0d",
        X"0404fb3d",
        X"0d780284",
        X"059f0533",
        X"70982b55",
        X"57557280",
        X"259b3875",
        X"80ff0656",
        X"805280f7",
        X"51e03f83",
        X"e0800881",
        X"ff065473",
        X"812680ff",
        X"388051fe",
        X"e73fffa2",
        X"3f8151fe",
        X"df3fff9a",
        X"3f7551fe",
        X"ed3f7498",
        X"2a51fee6",
        X"3f74902a",
        X"7081ff06",
        X"5253feda",
        X"3f74882a",
        X"7081ff06",
        X"5253fece",
        X"3f7481ff",
        X"0651fec6",
        X"3f815575",
        X"80c02e09",
        X"81068638",
        X"8195558d",
        X"397580c8",
        X"2e098106",
        X"84388187",
        X"557451fe",
        X"a53f8a55",
        X"fec83f83",
        X"e0800881",
        X"ff067098",
        X"2b545472",
        X"80258c38",
        X"ff157081",
        X"ff065653",
        X"74e23873",
        X"83e0800c",
        X"873d0d04",
        X"fa3d0dfd",
        X"c53f8051",
        X"fdda3f8a",
        X"54fe933f",
        X"ff147081",
        X"ff065553",
        X"73f33873",
        X"74535580",
        X"c051fea6",
        X"3f83e080",
        X"0881ff06",
        X"5473812e",
        X"09810682",
        X"a43883aa",
        X"5280c851",
        X"fe8c3f83",
        X"e0800881",
        X"ff065372",
        X"812e0981",
        X"0681ad38",
        X"7454883d",
        X"7405fc05",
        X"53fdc73f",
        X"83e08008",
        X"73348114",
        X"7081ff06",
        X"55538374",
        X"27e43802",
        X"9a053353",
        X"72812e09",
        X"810681dd",
        X"38029b05",
        X"335380ce",
        X"90547281",
        X"aa2e8d38",
        X"81cb3980",
        X"e4518ae0",
        X"3fff1454",
        X"73802e81",
        X"bc38820a",
        X"5281e951",
        X"fda43f83",
        X"e0800881",
        X"ff065372",
        X"de387252",
        X"80fa51fd",
        X"913f83e0",
        X"800881ff",
        X"06537281",
        X"94387254",
        X"883d7405",
        X"fc0553fc",
        X"d13f83e0",
        X"80087334",
        X"81147081",
        X"ff065553",
        X"837427e4",
        X"38873d33",
        X"70862a70",
        X"81065154",
        X"568c5572",
        X"80e33884",
        X"5580de39",
        X"745281e9",
        X"51fcc73f",
        X"83e08008",
        X"81ff0653",
        X"825581e9",
        X"56817327",
        X"86387355",
        X"80c15680",
        X"ce90548a",
        X"3980e451",
        X"89ce3fff",
        X"14547380",
        X"2ea93880",
        X"527551fc",
        X"953f83e0",
        X"800881ff",
        X"065372e1",
        X"38848052",
        X"80d051fc",
        X"813f83e0",
        X"800881ff",
        X"06537280",
        X"2e833880",
        X"557483e3",
        X"ac348051",
        X"fb823ffb",
        X"bd3f883d",
        X"0d04fb3d",
        X"0d775480",
        X"0b83e3ac",
        X"3370832a",
        X"70810651",
        X"55575572",
        X"752e0981",
        X"06853873",
        X"892b5473",
        X"5280d151",
        X"fbb83f83",
        X"e0800881",
        X"ff065372",
        X"bd3882b8",
        X"c054fafe",
        X"3f83e080",
        X"0881ff06",
        X"537281ff",
        X"2e098106",
        X"8938ff14",
        X"5473e738",
        X"9f397281",
        X"fe2e0981",
        X"06963883",
        X"e7b05283",
        X"e3b051fa",
        X"e83fface",
        X"3ffacb3f",
        X"83398155",
        X"8051fa84",
        X"3ffabf3f",
        X"7481ff06",
        X"83e0800c",
        X"873d0d04",
        X"fb3d0d77",
        X"83e3b056",
        X"548151f9",
        X"e73f83e3",
        X"ac337083",
        X"2a708106",
        X"51545672",
        X"85387389",
        X"2b547352",
        X"80d851fa",
        X"b13f83e0",
        X"800881ff",
        X"06537280",
        X"e43881ff",
        X"51f9cf3f",
        X"81fe51f9",
        X"c93f8480",
        X"53747081",
        X"05563351",
        X"f9bc3fff",
        X"137083ff",
        X"ff065153",
        X"72eb3872",
        X"51f9ab3f",
        X"7251f9a6",
        X"3ff9cb3f",
        X"83e08008",
        X"9f0653a7",
        X"88547285",
        X"2e8c3899",
        X"3980e451",
        X"87863fff",
        X"1454f9ae",
        X"3f83e080",
        X"0881ff2e",
        X"843873e9",
        X"388051f8",
        X"df3ff99a",
        X"3f800b83",
        X"e0800c87",
        X"3d0d0471",
        X"83e7b40c",
        X"8880800b",
        X"83e7b00c",
        X"8480800b",
        X"83e7b80c",
        X"04f13d0d",
        X"83808056",
        X"83e7b408",
        X"1683e7b0",
        X"08175654",
        X"74337434",
        X"83e7b808",
        X"16548074",
        X"34811656",
        X"758380a0",
        X"2e098106",
        X"db3883d0",
        X"805683e7",
        X"b4081683",
        X"e7b00817",
        X"56547433",
        X"743483e7",
        X"b8081654",
        X"80743481",
        X"16567583",
        X"d0902e09",
        X"8106db38",
        X"83a88056",
        X"83e7b408",
        X"1683e7b0",
        X"08175654",
        X"74337434",
        X"83e7b808",
        X"16548074",
        X"34811656",
        X"7583a890",
        X"2e098106",
        X"db388056",
        X"83e7b408",
        X"1683e7b8",
        X"08175555",
        X"73337534",
        X"81165675",
        X"8180802e",
        X"098106e4",
        X"3887ac3f",
        X"883d54a2",
        X"5380e8b8",
        X"5273519c",
        X"af3f8055",
        X"8c807458",
        X"5683e7b8",
        X"08165476",
        X"70810558",
        X"33743481",
        X"16811656",
        X"5674a22e",
        X"098106e5",
        X"38860b87",
        X"a8833480",
        X"0b87a882",
        X"34800b87",
        X"809a34af",
        X"0b878096",
        X"34bf0b87",
        X"80973480",
        X"0b878098",
        X"349f0b87",
        X"80993480",
        X"0b87809b",
        X"34f80b87",
        X"a8893474",
        X"87a88034",
        X"820b87d0",
        X"8f34820b",
        X"87a88134",
        X"840b8780",
        X"9f34ff0b",
        X"87d08b34",
        X"913d0d04",
        X"fe3d0d80",
        X"5383e7b8",
        X"081383e7",
        X"b4081452",
        X"52703372",
        X"34811353",
        X"72818080",
        X"2e098106",
        X"e4388380",
        X"805383e7",
        X"b8081383",
        X"e7b40814",
        X"52527033",
        X"72348113",
        X"53728380",
        X"a02e0981",
        X"06e43883",
        X"d0805383",
        X"e7b80813",
        X"83e7b408",
        X"14525270",
        X"33723481",
        X"13537283",
        X"d0902e09",
        X"8106e438",
        X"83a88053",
        X"83e7b808",
        X"1383e7b4",
        X"08145252",
        X"70337234",
        X"81135372",
        X"83a8902e",
        X"098106e4",
        X"38843d0d",
        X"04803d0d",
        X"90809008",
        X"810683e0",
        X"800c823d",
        X"0d04ff3d",
        X"0d908090",
        X"700870fe",
        X"06760772",
        X"0c525283",
        X"3d0d0480",
        X"3d0d9080",
        X"90087081",
        X"2c810683",
        X"e0800c51",
        X"823d0d04",
        X"ff3d0d90",
        X"80907008",
        X"70fd0676",
        X"1007720c",
        X"5252833d",
        X"0d04803d",
        X"0d908090",
        X"0870822c",
        X"bf0683e0",
        X"800c5182",
        X"3d0d04ff",
        X"3d0d9080",
        X"90700870",
        X"fe830676",
        X"822b0772",
        X"0c525283",
        X"3d0d0480",
        X"3d0d9080",
        X"90087088",
        X"2c870683",
        X"e0800c51",
        X"823d0d04",
        X"ff3d0d90",
        X"80907008",
        X"70f1ff06",
        X"76882b07",
        X"720c5252",
        X"833d0d04",
        X"803d0d90",
        X"80900870",
        X"912cbf06",
        X"83e0800c",
        X"51823d0d",
        X"04ff3d0d",
        X"90809070",
        X"0870fc87",
        X"ffff0676",
        X"912b0772",
        X"0c525283",
        X"3d0d0480",
        X"3d0d9080",
        X"90087099",
        X"2c810683",
        X"e0800c51",
        X"823d0d04",
        X"ff3d0d90",
        X"80907008",
        X"70ffbf0a",
        X"0676992b",
        X"07720c52",
        X"52833d0d",
        X"04803d0d",
        X"90808008",
        X"70882c81",
        X"0683e080",
        X"0c51823d",
        X"0d04803d",
        X"0d908080",
        X"0870892c",
        X"810683e0",
        X"800c5182",
        X"3d0d0480",
        X"3d0d9080",
        X"8008708a",
        X"2c810683",
        X"e0800c51",
        X"823d0d04",
        X"803d0d90",
        X"80800870",
        X"8b2c8106",
        X"83e0800c",
        X"51823d0d",
        X"04803d0d",
        X"90808008",
        X"70922c81",
        X"0683e080",
        X"0c51823d",
        X"0d04803d",
        X"0d908080",
        X"08708c2c",
        X"bf0683e0",
        X"800c5182",
        X"3d0d0480",
        X"3d0d9080",
        X"84088706",
        X"83e0800c",
        X"823d0d04",
        X"fe3d0d74",
        X"81e62987",
        X"2a9080a0",
        X"0c843d0d",
        X"04fe3d0d",
        X"7575ff19",
        X"53535370",
        X"ff2e8d38",
        X"72727081",
        X"055434ff",
        X"1151f039",
        X"843d0d04",
        X"fe3d0d75",
        X"75ff1953",
        X"535370ff",
        X"2e8d3872",
        X"72708405",
        X"540cff11",
        X"51f03984",
        X"3d0d04fe",
        X"3d0d8180",
        X"80538052",
        X"88800a51",
        X"ffb33fa0",
        X"80538052",
        X"82800a51",
        X"c73f843d",
        X"0d04803d",
        X"0d8151fc",
        X"853f7280",
        X"2e903880",
        X"51fdd93f",
        X"ce3f80eb",
        X"b83351fd",
        X"cf3f8151",
        X"fc963f80",
        X"51fc913f",
        X"8051fbe2",
        X"3f823d0d",
        X"04fd3d0d",
        X"75528054",
        X"80ff7225",
        X"8838810b",
        X"ff801353",
        X"54ffbf12",
        X"51709926",
        X"8638e012",
        X"52b039ff",
        X"9f125199",
        X"7127a738",
        X"d012e013",
        X"54517089",
        X"26853872",
        X"52983972",
        X"8f268538",
        X"72528f39",
        X"71ba2e09",
        X"81068538",
        X"9a528339",
        X"80527380",
        X"2e853881",
        X"80125271",
        X"81ff0683",
        X"e0800c85",
        X"3d0d0480",
        X"3d0d84d8",
        X"c0518071",
        X"70810553",
        X"347084e0",
        X"c02e0981",
        X"06f03882",
        X"3d0d04fe",
        X"3d0d0297",
        X"053351fe",
        X"f43f83e0",
        X"800881ff",
        X"0683e7c0",
        X"08545280",
        X"73249b38",
        X"83e7e808",
        X"137283e7",
        X"ec080753",
        X"53717334",
        X"83e7c008",
        X"810583e7",
        X"c00c843d",
        X"0d04fa3d",
        X"0d82800a",
        X"1b558057",
        X"883dfc05",
        X"54795374",
        X"527851ff",
        X"b9d73f88",
        X"3d0d04fe",
        X"3d0d83e7",
        X"d8085274",
        X"51c0bb3f",
        X"83e08008",
        X"8c387653",
        X"755283e7",
        X"d80851c6",
        X"3f843d0d",
        X"04fe3d0d",
        X"83e7d808",
        X"53755274",
        X"51ffbaf9",
        X"3f83e080",
        X"088d3877",
        X"53765283",
        X"e7d80851",
        X"ffa03f84",
        X"3d0d04fd",
        X"3d0d83e7",
        X"d80851ff",
        X"b9ec3f83",
        X"e0800890",
        X"802e0981",
        X"06ad3880",
        X"5483c180",
        X"805383e0",
        X"80085283",
        X"e7d80851",
        X"fef03f87",
        X"c1808014",
        X"3387c190",
        X"80153481",
        X"14547390",
        X"802e0981",
        X"06e93885",
        X"3d0d04fc",
        X"3d0d7654",
        X"73902e80",
        X"ff387390",
        X"248e3873",
        X"842e9838",
        X"73862ea6",
        X"3882b939",
        X"73932e81",
        X"95387394",
        X"2e81cf38",
        X"82aa3981",
        X"80805382",
        X"80805283",
        X"e7d40851",
        X"fe983f82",
        X"b5398054",
        X"81808053",
        X"80c08052",
        X"83e7d408",
        X"51fe833f",
        X"82808053",
        X"80c08052",
        X"83e7d408",
        X"51fdf33f",
        X"84818080",
        X"14338481",
        X"c0801534",
        X"84828080",
        X"14338482",
        X"c0801534",
        X"81145473",
        X"80c0802e",
        X"098106dc",
        X"3881eb39",
        X"82808053",
        X"81808052",
        X"83e7d408",
        X"51fdbb3f",
        X"80548482",
        X"80801433",
        X"84818080",
        X"15348114",
        X"54738180",
        X"802e0981",
        X"06e83881",
        X"bd398180",
        X"805380c0",
        X"805283e7",
        X"d40851fd",
        X"8d3f8055",
        X"84818080",
        X"15547333",
        X"8481c080",
        X"16347333",
        X"84828080",
        X"16347333",
        X"8482c080",
        X"16348115",
        X"557480c0",
        X"802e0981",
        X"06d63880",
        X"fd398180",
        X"8053a080",
        X"5283e7d4",
        X"0851fcce",
        X"3f805584",
        X"81808015",
        X"54733384",
        X"81a08016",
        X"34733384",
        X"81c08016",
        X"34733384",
        X"81e08016",
        X"34733384",
        X"82808016",
        X"34733384",
        X"82a08016",
        X"34733384",
        X"82c08016",
        X"34733384",
        X"82e08016",
        X"34811555",
        X"74a0802e",
        X"098106ff",
        X"b6389f39",
        X"fba53f80",
        X"0b83e7c0",
        X"0c800b83",
        X"e7ec0c80",
        X"e99c51e7",
        X"d83f81b7",
        X"8dc051f9",
        X"873f863d",
        X"0d04fc3d",
        X"0d767052",
        X"55ffbd96",
        X"3f83e080",
        X"08548153",
        X"83e08008",
        X"80c23874",
        X"51ffbcd8",
        X"3f83e080",
        X"0880e9b8",
        X"5383e080",
        X"085253d5",
        X"b63f83e0",
        X"8008a138",
        X"80e9bc52",
        X"7251d5a7",
        X"3f83e080",
        X"08923880",
        X"e9c05272",
        X"51d5983f",
        X"83e08008",
        X"802e8338",
        X"81547353",
        X"7283e080",
        X"0c863d0d",
        X"04f13d0d",
        X"80d6e20b",
        X"83e3900c",
        X"83e7d408",
        X"51d7b63f",
        X"83e08008",
        X"5583e080",
        X"08802e81",
        X"ea3883e7",
        X"d40851ff",
        X"b2af3fff",
        X"0b80e9bc",
        X"5383e080",
        X"085256d4",
        X"ca3f83e0",
        X"8008802e",
        X"9f388058",
        X"913ddc11",
        X"55559053",
        X"f0155283",
        X"e7d40851",
        X"ffb4923f",
        X"02b70533",
        X"5681a539",
        X"83e7d408",
        X"51ffb4ee",
        X"3f83e080",
        X"085783e0",
        X"80088280",
        X"802e0981",
        X"06833884",
        X"5683e080",
        X"08818080",
        X"2e098106",
        X"80e13880",
        X"5c805b80",
        X"5a8059f9",
        X"8e3f800b",
        X"83e7c00c",
        X"800b83e7",
        X"ec0c80e9",
        X"c451e5c1",
        X"3f80d00b",
        X"83e7c00c",
        X"80e9d451",
        X"e5b33f80",
        X"f80b83e7",
        X"c00c80e9",
        X"e851e5a5",
        X"3f758025",
        X"a2388052",
        X"893d7052",
        X"558ad73f",
        X"83527451",
        X"8ad03f78",
        X"55748025",
        X"83389056",
        X"807525dd",
        X"38865676",
        X"80c0802e",
        X"09810685",
        X"3893568c",
        X"3976a080",
        X"2e098106",
        X"83389456",
        X"7551fa9f",
        X"3f815574",
        X"83e0800c",
        X"913d0d04",
        X"f73d0d80",
        X"5a805980",
        X"58805780",
        X"705656f7",
        X"fe3f800b",
        X"83e7c00c",
        X"800b83e7",
        X"ec0c80e9",
        X"fc51e4b1",
        X"3f81800b",
        X"83e7ec0c",
        X"80ea8051",
        X"e4a33f80",
        X"f80b83e7",
        X"c00c7430",
        X"70760780",
        X"2570872b",
        X"83e7ec0c",
        X"515383e7",
        X"d80851ff",
        X"aff33f83",
        X"e0800852",
        X"80ea8851",
        X"e3f73f81",
        X"c80b83e7",
        X"c00c7481",
        X"32703070",
        X"72078025",
        X"70872b83",
        X"e7ec0c51",
        X"5483e7d4",
        X"085254ff",
        X"afc33f80",
        X"ea905383",
        X"e0800880",
        X"2e8f3883",
        X"e7d40851",
        X"ffafae3f",
        X"83e08008",
        X"53725280",
        X"ea9851e3",
        X"b03f82c0",
        X"0b83e7c0",
        X"0c748232",
        X"70307072",
        X"07802570",
        X"872b83e7",
        X"ec0c5154",
        X"80eaa052",
        X"54e38e3f",
        X"868da051",
        X"f4be3ff3",
        X"eb3f83e0",
        X"8008f838",
        X"83e08008",
        X"52873d70",
        X"525388b2",
        X"3f835272",
        X"5188ab3f",
        X"79537280",
        X"ef387715",
        X"55748025",
        X"86388255",
        X"80d93982",
        X"75258538",
        X"72559a39",
        X"74812eb9",
        X"38748124",
        X"89387480",
        X"2e8b3880",
        X"c1397482",
        X"2eb938ba",
        X"39768638",
        X"78802eb2",
        X"3883e38c",
        X"0883e388",
        X"0caedb0b",
        X"83e3900c",
        X"83e7d808",
        X"51d2f63f",
        X"f7893f96",
        X"39768638",
        X"78802e8e",
        X"38fb9e3f",
        X"83e08008",
        X"538c3978",
        X"87387580",
        X"2efdb038",
        X"80537283",
        X"e0800c8b",
        X"3d0d04f9",
        X"3d0d8058",
        X"80578056",
        X"8055f285",
        X"3f83e080",
        X"08802e86",
        X"38805181",
        X"8a39f28a",
        X"3f83e080",
        X"0880fe38",
        X"f2aa3f83",
        X"e0800880",
        X"2ebd3881",
        X"51efe73f",
        X"ec9f3f80",
        X"0b83e7c0",
        X"0cfcd53f",
        X"83e08008",
        X"53805289",
        X"3df00551",
        X"86dc3ff1",
        X"ff3f83e0",
        X"8008f838",
        X"ff0b83e7",
        X"c00ceea0",
        X"3f72be38",
        X"7251efb2",
        X"3fbc39f1",
        X"ce3f83e0",
        X"8008802e",
        X"b1388151",
        X"efa03feb",
        X"d83ffa81",
        X"3f83e080",
        X"08538052",
        X"893df005",
        X"51869b3f",
        X"f1be3f83",
        X"e08008f8",
        X"38ede53f",
        X"72802e86",
        X"388151f2",
        X"e93f893d",
        X"0d04fe3d",
        X"0d828080",
        X"53805281",
        X"81808051",
        X"f1f73f80",
        X"c0805380",
        X"52848180",
        X"8051f288",
        X"3f908080",
        X"52868480",
        X"8051ffb0",
        X"aa3f83e0",
        X"8008a438",
        X"80ebbc51",
        X"ffb4ed3f",
        X"83e7d808",
        X"5380eaa8",
        X"5283e080",
        X"0851ffaf",
        X"cc3f83e0",
        X"80088438",
        X"f4e13f81",
        X"51f28b3f",
        X"fdf93ffc",
        X"3983e08c",
        X"080283e0",
        X"8c0cfb3d",
        X"0d0280ea",
        X"b40b83e3",
        X"8c0c80e9",
        X"c00b83e3",
        X"840c80e9",
        X"bc0b83e3",
        X"980c80ea",
        X"b80b83e3",
        X"940c83e0",
        X"8c08fc05",
        X"0c800b83",
        X"e7c40b83",
        X"e08c08f8",
        X"050c83e0",
        X"8c08f405",
        X"0cffaea3",
        X"3f83e080",
        X"088605fc",
        X"0683e08c",
        X"08f0050c",
        X"0283e08c",
        X"08f00508",
        X"310d833d",
        X"7083e08c",
        X"08f80508",
        X"70840583",
        X"e08c08f8",
        X"050c0c51",
        X"ffaae43f",
        X"83e08c08",
        X"f4050881",
        X"0583e08c",
        X"08f4050c",
        X"83e08c08",
        X"f4050889",
        X"2e098106",
        X"ffab3886",
        X"94808051",
        X"e9913fff",
        X"0b83e7c0",
        X"0c800b83",
        X"e7ec0c84",
        X"d8c00b83",
        X"e7e80c81",
        X"51ecd33f",
        X"8151ecf8",
        X"3f8051ec",
        X"f33fed86",
        X"3f83e080",
        X"088b3881",
        X"51ed903f",
        X"8251edb8",
        X"3f8051ed",
        X"e03f8051",
        X"ee8a3f80",
        X"d2835280",
        X"51dde73f",
        X"fdb03f83",
        X"e08c08fc",
        X"05080d80",
        X"0b83e080",
        X"0c873d0d",
        X"83e08c0c",
        X"04fb3d0d",
        X"77548074",
        X"0c800b84",
        X"150c800b",
        X"88150c80",
        X"0b8c150c",
        X"eed03f83",
        X"e0800887",
        X"d0883370",
        X"81ff0651",
        X"525570a7",
        X"3887d080",
        X"3383e7fc",
        X"3487d081",
        X"3383e7f8",
        X"3487d082",
        X"3383e7f0",
        X"3487d083",
        X"3383e7f4",
        X"34ff0b87",
        X"d08b3487",
        X"d0893387",
        X"d08f3370",
        X"822a7081",
        X"06703070",
        X"72077009",
        X"709f2c77",
        X"069e0657",
        X"51515551",
        X"51535380",
        X"73980652",
        X"5270882e",
        X"09810683",
        X"38815270",
        X"98327030",
        X"70802574",
        X"71318418",
        X"0c515151",
        X"80738606",
        X"52527082",
        X"2e098106",
        X"83388152",
        X"70863270",
        X"30708025",
        X"74713177",
        X"0c515151",
        X"83e7fc33",
        X"5181aa71",
        X"27843881",
        X"740c83e7",
        X"fc335170",
        X"bb268438",
        X"ff740c83",
        X"e7f83351",
        X"81aa7127",
        X"8638810b",
        X"84150c83",
        X"e7f83351",
        X"70bb2686",
        X"38ff0b84",
        X"150c83e7",
        X"f0335181",
        X"aa712784",
        X"3881740c",
        X"83e7f033",
        X"5170bb26",
        X"8438ff74",
        X"0c83e7f4",
        X"335181aa",
        X"71278638",
        X"810b8415",
        X"0c83e7f4",
        X"335170bb",
        X"268638ff",
        X"0b84150c",
        X"80567294",
        X"2eaa3887",
        X"80903387",
        X"80913387",
        X"80923370",
        X"81ff0672",
        X"74060687",
        X"80933371",
        X"06810651",
        X"52535353",
        X"71762e09",
        X"81068338",
        X"81567588",
        X"150c7480",
        X"2eb03874",
        X"812a7081",
        X"06768106",
        X"3184160c",
        X"5174832a",
        X"75822a71",
        X"81067181",
        X"0631760c",
        X"52527484",
        X"2a810688",
        X"150c7485",
        X"2a81068c",
        X"150c873d",
        X"0d04fe3d",
        X"0d747654",
        X"527151fc",
        X"dc3feb98",
        X"3f83e080",
        X"08802e89",
        X"38810b8c",
        X"130c80d0",
        X"3972812e",
        X"a7388173",
        X"268d3872",
        X"822ead38",
        X"72832ea1",
        X"38d33971",
        X"08cf3884",
        X"1208ca38",
        X"881208c5",
        X"388c1208",
        X"c038a539",
        X"88120881",
        X"2e9e3891",
        X"39881208",
        X"812e9538",
        X"71089138",
        X"8412088c",
        X"388c1208",
        X"812e0981",
        X"06ff9a38",
        X"843d0d04",
        X"fe3d0d80",
        X"53755274",
        X"5181923f",
        X"843d0d04",
        X"fe3d0d81",
        X"53755274",
        X"5181823f",
        X"843d0d04",
        X"fb3d0d77",
        X"79555580",
        X"56747625",
        X"86387430",
        X"55815673",
        X"80258838",
        X"73307681",
        X"32575480",
        X"53735274",
        X"5180d63f",
        X"83e08008",
        X"5475802e",
        X"873883e0",
        X"80083054",
        X"7383e080",
        X"0c873d0d",
        X"04fa3d0d",
        X"787a5755",
        X"80577477",
        X"25863874",
        X"30558157",
        X"759f2c54",
        X"81537574",
        X"32743152",
        X"74519a3f",
        X"83e08008",
        X"5476802e",
        X"873883e0",
        X"80083054",
        X"7383e080",
        X"0c883d0d",
        X"04fc3d0d",
        X"76785354",
        X"81538055",
        X"87397110",
        X"73105452",
        X"73722651",
        X"72802ea7",
        X"3870802e",
        X"86387180",
        X"25e83872",
        X"802e9838",
        X"71742689",
        X"38737231",
        X"75740756",
        X"5472812a",
        X"72812a53",
        X"53e53973",
        X"51788338",
        X"74517083",
        X"e0800c86",
        X"3d0d04fd",
        X"3d0d7577",
        X"54528054",
        X"718106ff",
        X"11700975",
        X"06167481",
        X"2a761057",
        X"55565151",
        X"71ea3873",
        X"83e0800c",
        X"853d0d04",
        X"fd3d0d75",
        X"7771ff1b",
        X"54565452",
        X"70ff2e92",
        X"38727081",
        X"05543372",
        X"70810554",
        X"34ff1151",
        X"eb397383",
        X"e0800c85",
        X"3d0d0400",
        X"00ffffff",
        X"ff00ffff",
        X"ffff00ff",
        X"ffffff00",
        X"809a9041",
        X"8e418f80",
        X"45454549",
        X"49498e8f",
        X"9092924f",
        X"994f5555",
        X"59999a9b",
        X"9c9d9e9f",
        X"41494f55",
        X"a5a5a6a7",
        X"a8a9aaab",
        X"ac21aeaf",
        X"b0b1b2b3",
        X"b4b5b6b7",
        X"b8b9babb",
        X"bcbdbebf",
        X"c0c1c2c3",
        X"c4c5c6c7",
        X"c8c9cacb",
        X"cccdcecf",
        X"d0d1d2d3",
        X"d4d5d6d7",
        X"d8d9dadb",
        X"dcdddedf",
        X"e0e1e2e3",
        X"e4e5e6e7",
        X"e8e9eaeb",
        X"ecedeeef",
        X"f0f1f2f3",
        X"f4f5f6f7",
        X"f8f9fafb",
        X"fcfdfeff",
        X"00000000",
        X"70704740",
        X"2c704268",
        X"2c020202",
        X"02020202",
        X"02020202",
        X"02020202",
        X"02020202",
        X"02020241",
        X"00060000",
        X"2e2e0000",
        X"41545200",
        X"58464400",
        X"58455800",
        X"43686f6f",
        X"73652000",
        X"66696c65",
        X"00000000",
        X"4449523a",
        X"00000000",
        X"44495200",
        X"25732025",
        X"73000000",
        X"20000000",
        X"25303278",
        X"00000000",
        X"556e6b6e",
        X"6f776e20",
        X"74797065",
        X"206f6620",
        X"63617274",
        X"72696467",
        X"65210000",
        X"41353200",
        X"43415200",
        X"42494e00",
        X"31366b20",
        X"63617274",
        X"20747970",
        X"65000000",
        X"4c656674",
        X"20666f72",
        X"206f6e65",
        X"20636869",
        X"70000000",
        X"52696768",
        X"7420666f",
        X"72207477",
        X"6f206368",
        X"69700000",
        X"53650000",
        X"7474696e",
        X"67730000",
        X"526f6d3a",
        X"25730000",
        X"4e4f4e45",
        X"00000000",
        X"43617274",
        X"3a257300",
        X"45786974",
        X"00000000",
        X"35323030",
        X"2e726f6d",
        X"00000000",
        X"524f4d00",
        X"4d454d00",
        X"00000000",
        X"00000000",
        X"01010008",
        X"02210010",
        X"080d0040",
        X"090a0040",
        X"0a090040",
        X"0b080040",
        X"0c300020",
        X"0d310040",
        X"0e320080",
        X"0f040010",
        X"110c0080",
        X"17330100",
        X"18340200",
        X"1a280010",
        X"1b290020",
        X"1c2a0040",
        X"1d2b0080",
        X"1e2c0100",
        X"1f2d0200",
        X"21380020",
        X"22390040",
        X"233a0080",
        X"243b0100",
        X"253c0200",
        X"28230010",
        X"29020080",
        X"2a030400",
        X"38240200",
        X"00000000",
        X"00000000",
        X"2f617461",
        X"72353230",
        X"302f726f",
        X"6d000000",
        X"2f617461",
        X"72353230",
        X"302f7573",
        X"65720000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000"

);

signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
