
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(12 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 8191) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
        X"0b0b0b89",
        X"ad040b0b",
        X"0b0b0b0b",
        X"0b0b0b0b",
        X"0b0b0b0b",
        X"0b0b0b0b",
        X"0b0b0b0b",
        X"0b0b0b0b",
        X"0b0b0b0b",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"71fd0608",
        X"72830609",
        X"81058205",
        X"832b2a83",
        X"ffff0652",
        X"04000000",
        X"00000000",
        X"00000000",
        X"71fd0608",
        X"83ffff73",
        X"83060981",
        X"05820583",
        X"2b2b0906",
        X"7383ffff",
        X"0b0b0b0b",
        X"83a70400",
        X"72098105",
        X"72057373",
        X"09060906",
        X"73097306",
        X"070a8106",
        X"53510400",
        X"00000000",
        X"00000000",
        X"72722473",
        X"732e0753",
        X"51040000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"71737109",
        X"71068106",
        X"30720a10",
        X"0a720a10",
        X"0a31050a",
        X"81065151",
        X"53510400",
        X"00000000",
        X"72722673",
        X"732e0753",
        X"51040000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"0b0b0b88",
        X"bc040000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"720a722b",
        X"0a535104",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"72729f06",
        X"0981050b",
        X"0b0b889f",
        X"05040000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"72722aff",
        X"739f062a",
        X"0974090a",
        X"8106ff05",
        X"06075351",
        X"04000000",
        X"00000000",
        X"00000000",
        X"71715351",
        X"020d0406",
        X"73830609",
        X"81058205",
        X"832b0b2b",
        X"0772fc06",
        X"0c515104",
        X"00000000",
        X"72098105",
        X"72050970",
        X"81050906",
        X"0a810653",
        X"51040000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"72098105",
        X"72050970",
        X"81050906",
        X"0a098106",
        X"53510400",
        X"00000000",
        X"00000000",
        X"00000000",
        X"71098105",
        X"52040000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"72720981",
        X"05055351",
        X"04000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"72097206",
        X"73730906",
        X"07535104",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"71fc0608",
        X"72830609",
        X"81058305",
        X"1010102a",
        X"81ff0652",
        X"04000000",
        X"00000000",
        X"00000000",
        X"71fc0608",
        X"0b0b80f8",
        X"f0738306",
        X"10100508",
        X"060b0b0b",
        X"88a20400",
        X"00000000",
        X"00000000",
        X"0b0b0b88",
        X"ff040000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"0b0b0b88",
        X"d8040000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"72097081",
        X"0509060a",
        X"8106ff05",
        X"70547106",
        X"73097274",
        X"05ff0506",
        X"07515151",
        X"04000000",
        X"72097081",
        X"0509060a",
        X"098106ff",
        X"05705471",
        X"06730972",
        X"7405ff05",
        X"06075151",
        X"51040000",
        X"05ff0504",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"810b80fc",
        X"ac0c5104",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00007181",
        X"05520400",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000284",
        X"05721010",
        X"05520400",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00007171",
        X"05ff0571",
        X"5351020d",
        X"04000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"10101010",
        X"10101010",
        X"10101010",
        X"10101010",
        X"10101010",
        X"10101010",
        X"10101010",
        X"10101053",
        X"51047381",
        X"ff067383",
        X"06098105",
        X"83051010",
        X"102b0772",
        X"fc060c51",
        X"51043c04",
        X"72728072",
        X"8106ff05",
        X"09720605",
        X"71105272",
        X"0a100a53",
        X"72ed3851",
        X"51535104",
        X"83c08008",
        X"83c08408",
        X"83c08808",
        X"757580f6",
        X"842d5050",
        X"83c08008",
        X"5683c088",
        X"0c83c084",
        X"0c83c080",
        X"0c510483",
        X"c0800883",
        X"c0840883",
        X"c0880875",
        X"7580f5c3",
        X"2d505083",
        X"c0800856",
        X"83c0880c",
        X"83c0840c",
        X"83c0800c",
        X"51040000",
        X"800489aa",
        X"0489aa0b",
        X"80dfa104",
        X"fd3d0d75",
        X"705254af",
        X"be3f83c0",
        X"80081453",
        X"72742e92",
        X"38ff1370",
        X"33535371",
        X"af2e0981",
        X"06ee3881",
        X"13537283",
        X"c0800c85",
        X"3d0d04fd",
        X"3d0d7577",
        X"70535454",
        X"c73f83c0",
        X"8008732e",
        X"a13883c0",
        X"80087331",
        X"52ff1252",
        X"71ff2e8f",
        X"38727081",
        X"05543374",
        X"70810556",
        X"34eb39ff",
        X"14548074",
        X"34853d0d",
        X"04803d0d",
        X"7251ff90",
        X"3f823d0d",
        X"047183c0",
        X"800c0480",
        X"3d0d7251",
        X"80713481",
        X"0bbc120c",
        X"800b80c0",
        X"120c823d",
        X"0d04800b",
        X"83c2c408",
        X"248a38b6",
        X"8f3fff0b",
        X"83c2c40c",
        X"800b83c0",
        X"800c04ff",
        X"3d0d7352",
        X"83c0a008",
        X"722e8d38",
        X"d93f7151",
        X"96a03f71",
        X"83c0a00c",
        X"833d0d04",
        X"f43d0d7e",
        X"60625c5a",
        X"55805681",
        X"54bc1508",
        X"762e0981",
        X"06819138",
        X"7451c83f",
        X"7958757a",
        X"2580f738",
        X"83c2f408",
        X"70892a57",
        X"83ff0678",
        X"84807231",
        X"56565773",
        X"78258338",
        X"73557583",
        X"c2c4082e",
        X"8438ff82",
        X"3f83c2c4",
        X"088025a6",
        X"3875892b",
        X"5198dc3f",
        X"83c2f408",
        X"8f3dfc11",
        X"555c5481",
        X"52f81b51",
        X"96c63f76",
        X"1483c2f4",
        X"0c7583c2",
        X"c40c7453",
        X"76527851",
        X"b4b93f83",
        X"c0800883",
        X"c2f40816",
        X"83c2f40c",
        X"78763176",
        X"1b5b5956",
        X"778024ff",
        X"8b38617a",
        X"710c5475",
        X"5475802e",
        X"83388154",
        X"7383c080",
        X"0c8e3d0d",
        X"04fc3d0d",
        X"fe943f76",
        X"51fea83f",
        X"863dfc05",
        X"53785277",
        X"5195e93f",
        X"7975710c",
        X"5483c080",
        X"085483c0",
        X"8008802e",
        X"83388154",
        X"7383c080",
        X"0c863d0d",
        X"04fe3d0d",
        X"7583c2c4",
        X"08535380",
        X"72248938",
        X"71732e84",
        X"38fdcf3f",
        X"7451fde3",
        X"3f725197",
        X"ae3f83c0",
        X"80085283",
        X"c0800880",
        X"2e833881",
        X"527183c0",
        X"800c843d",
        X"0d04803d",
        X"0d7280c0",
        X"110883c0",
        X"800c5182",
        X"3d0d0480",
        X"3d0d72bc",
        X"110883c0",
        X"800c5182",
        X"3d0d0480",
        X"c40b83c0",
        X"800c04fd",
        X"3d0d7577",
        X"71547053",
        X"5553ab8f",
        X"3f82c813",
        X"08bc150c",
        X"82c01308",
        X"80c0150c",
        X"fce43f73",
        X"5193ab3f",
        X"7383c0a0",
        X"0c83c080",
        X"085383c0",
        X"8008802e",
        X"83388153",
        X"7283c080",
        X"0c853d0d",
        X"04fd3d0d",
        X"75775553",
        X"fcb83f72",
        X"802ea538",
        X"bc130852",
        X"7351aa99",
        X"3f83c080",
        X"088f3877",
        X"527251ff",
        X"9a3f83c0",
        X"8008538a",
        X"3982cc13",
        X"0853d839",
        X"81537283",
        X"c0800c85",
        X"3d0d04fe",
        X"3d0dff0b",
        X"83c2c40c",
        X"7483c0a4",
        X"0c7583c2",
        X"c00cb0ed",
        X"3f83c080",
        X"0881ff06",
        X"52815371",
        X"993883c2",
        X"dc518e94",
        X"3f83c080",
        X"085283c0",
        X"8008802e",
        X"83387252",
        X"71537283",
        X"c0800c84",
        X"3d0d04fa",
        X"3d0d787a",
        X"82c41208",
        X"82c41208",
        X"70722459",
        X"56565757",
        X"73732e09",
        X"81069138",
        X"80c01652",
        X"80c01751",
        X"a88a3f83",
        X"c0800855",
        X"7483c080",
        X"0c883d0d",
        X"04f63d0d",
        X"7c5b807b",
        X"715c5457",
        X"7a772e8c",
        X"38811a82",
        X"cc140854",
        X"5a72f638",
        X"805980d9",
        X"397a5481",
        X"5780707b",
        X"7b315a57",
        X"55ff1853",
        X"74732580",
        X"c13882cc",
        X"14085273",
        X"51ff8c3f",
        X"800b83c0",
        X"800825a1",
        X"3882cc14",
        X"0882cc11",
        X"0882cc16",
        X"0c7482cc",
        X"120c5375",
        X"802e8638",
        X"7282cc17",
        X"0c725480",
        X"577382cc",
        X"15088117",
        X"575556ff",
        X"b8398119",
        X"59800bff",
        X"1b545478",
        X"73258338",
        X"81547681",
        X"32707506",
        X"515372ff",
        X"90388c3d",
        X"0d04f73d",
        X"0d7b7d5a",
        X"5a82d052",
        X"83c2c008",
        X"5180e4bf",
        X"3f83c080",
        X"0857f9da",
        X"3f795283",
        X"c2c85195",
        X"b73f83c0",
        X"80085480",
        X"5383c080",
        X"08732e09",
        X"81068283",
        X"3883c0a4",
        X"080b0b80",
        X"faa05370",
        X"5256a7c7",
        X"3f0b0b80",
        X"faa05280",
        X"c01651a7",
        X"ba3f75bc",
        X"170c7382",
        X"c0170c81",
        X"0b82c417",
        X"0c810b82",
        X"c8170c73",
        X"82cc170c",
        X"ff1782d0",
        X"17555781",
        X"913983c0",
        X"b0337082",
        X"2a708106",
        X"51545572",
        X"81803874",
        X"812a8106",
        X"587780f6",
        X"3874842a",
        X"810682c4",
        X"150c83c0",
        X"b0338106",
        X"82c8150c",
        X"79527351",
        X"a6e13f73",
        X"51a6f83f",
        X"83c08008",
        X"1453af73",
        X"70810555",
        X"3472bc15",
        X"0c83c0b1",
        X"527251a6",
        X"c23f83c0",
        X"a80882c0",
        X"150c83c0",
        X"be5280c0",
        X"1451a6af",
        X"3f78802e",
        X"8d387351",
        X"782d83c0",
        X"8008802e",
        X"99387782",
        X"cc150c75",
        X"802e8638",
        X"7382cc17",
        X"0c7382d0",
        X"15ff1959",
        X"55567680",
        X"2e9b3883",
        X"c0a85283",
        X"c2c85194",
        X"ad3f83c0",
        X"80088a38",
        X"83c0b133",
        X"5372fed2",
        X"3878802e",
        X"893883c0",
        X"a40851fc",
        X"b83f83c0",
        X"a4085372",
        X"83c0800c",
        X"8b3d0d04",
        X"ff3d0d80",
        X"527351fd",
        X"b53f833d",
        X"0d04f03d",
        X"0d627052",
        X"54f6893f",
        X"83c08008",
        X"7453873d",
        X"70535555",
        X"f6a93ff7",
        X"893f7351",
        X"d33f6353",
        X"745283c0",
        X"800851fa",
        X"b83f923d",
        X"0d047183",
        X"c0800c04",
        X"80c01283",
        X"c0800c04",
        X"803d0d72",
        X"82c01108",
        X"83c0800c",
        X"51823d0d",
        X"04803d0d",
        X"7282cc11",
        X"0883c080",
        X"0c51823d",
        X"0d04803d",
        X"0d7282c4",
        X"110883c0",
        X"800c5182",
        X"3d0d04f9",
        X"3d0d7983",
        X"c0900857",
        X"57817727",
        X"81963876",
        X"88170827",
        X"818e3875",
        X"33557482",
        X"2e893874",
        X"832eb338",
        X"80fe3974",
        X"54761083",
        X"fe065376",
        X"882a8c17",
        X"08055289",
        X"3dfc0551",
        X"ab9b3f83",
        X"c0800880",
        X"df38029d",
        X"0533893d",
        X"3371882b",
        X"07565680",
        X"d1398454",
        X"76822b83",
        X"fc065376",
        X"872a8c17",
        X"08055289",
        X"3dfc0551",
        X"aaeb3f83",
        X"c08008b0",
        X"38029f05",
        X"33028405",
        X"9e053371",
        X"982b7190",
        X"2b07028c",
        X"059d0533",
        X"70882b72",
        X"078d3d33",
        X"7180ffff",
        X"fe800607",
        X"51525357",
        X"58568339",
        X"81557483",
        X"c0800c89",
        X"3d0d04fb",
        X"3d0d83c0",
        X"9008fe19",
        X"881208fe",
        X"05555654",
        X"80567473",
        X"278d3882",
        X"14337571",
        X"29941608",
        X"05575375",
        X"83c0800c",
        X"873d0d04",
        X"fc3d0d76",
        X"52800b83",
        X"c0900870",
        X"33515253",
        X"70832e09",
        X"81069138",
        X"95123394",
        X"13337198",
        X"2b71902b",
        X"07555551",
        X"9b12339a",
        X"13337188",
        X"2b077407",
        X"83c0800c",
        X"55863d0d",
        X"04fc3d0d",
        X"7683c090",
        X"08555580",
        X"75238815",
        X"08537281",
        X"2e883888",
        X"14087326",
        X"85388152",
        X"b2397290",
        X"38733352",
        X"71832e09",
        X"81068538",
        X"90140853",
        X"728c160c",
        X"72802e8d",
        X"387251fe",
        X"d63f83c0",
        X"80085285",
        X"39901408",
        X"52719016",
        X"0c805271",
        X"83c0800c",
        X"863d0d04",
        X"fa3d0d78",
        X"83c09008",
        X"71228105",
        X"7083ffff",
        X"06575457",
        X"5573802e",
        X"88389015",
        X"08537286",
        X"38835280",
        X"e739738f",
        X"06527180",
        X"da388113",
        X"90160c8c",
        X"15085372",
        X"9038830b",
        X"84172257",
        X"52737627",
        X"80c638bf",
        X"39821633",
        X"ff057484",
        X"2a065271",
        X"b2387251",
        X"fcb13f81",
        X"527183c0",
        X"800827a8",
        X"38835283",
        X"c0800888",
        X"1708279c",
        X"3883c080",
        X"088c160c",
        X"83c08008",
        X"51fdbc3f",
        X"83c08008",
        X"90160c73",
        X"75238052",
        X"7183c080",
        X"0c883d0d",
        X"04f23d0d",
        X"60626458",
        X"5e5b7533",
        X"5574a02e",
        X"09810688",
        X"38811670",
        X"4456ef39",
        X"62703356",
        X"5674af2e",
        X"09810684",
        X"38811643",
        X"800b881c",
        X"0c627033",
        X"5155749f",
        X"2691387a",
        X"51fdd23f",
        X"83c08008",
        X"56807d34",
        X"83813993",
        X"3d841c08",
        X"7058595f",
        X"8a55a076",
        X"70810558",
        X"34ff1555",
        X"74ff2e09",
        X"8106ef38",
        X"80705a5c",
        X"887f085f",
        X"5a7b811d",
        X"7081ff06",
        X"60137033",
        X"70af3270",
        X"30a07327",
        X"71802507",
        X"5151525b",
        X"535e5755",
        X"7480e738",
        X"76ae2e09",
        X"81068338",
        X"8155787a",
        X"27750755",
        X"74802e9f",
        X"38798832",
        X"703078ae",
        X"32703070",
        X"73079f2a",
        X"53515751",
        X"5675bb38",
        X"88598b5a",
        X"ffab3976",
        X"982b5574",
        X"80258738",
        X"80f88017",
        X"3357ff9f",
        X"17557499",
        X"268938e0",
        X"177081ff",
        X"06585578",
        X"811a7081",
        X"ff067a13",
        X"535b5755",
        X"767534fe",
        X"f8397b1e",
        X"7f0c8055",
        X"76a02683",
        X"38815574",
        X"8b19347a",
        X"51fc823f",
        X"83c08008",
        X"80f538a0",
        X"547a2270",
        X"852b83e0",
        X"06545590",
        X"1b08527c",
        X"51a5a63f",
        X"83c08008",
        X"5783c080",
        X"08818138",
        X"7c335574",
        X"802e80f4",
        X"388b1d33",
        X"70832a70",
        X"81065156",
        X"5674b438",
        X"8b7d841d",
        X"0883c080",
        X"08595b5b",
        X"58ff1858",
        X"77ff2e9a",
        X"38797081",
        X"055b3379",
        X"7081055b",
        X"33717131",
        X"52565675",
        X"802ee238",
        X"86397580",
        X"2e96387a",
        X"51fbe53f",
        X"ff863983",
        X"c0800856",
        X"83c08008",
        X"b6388339",
        X"7656841b",
        X"088b1133",
        X"515574a7",
        X"388b1d33",
        X"70842a70",
        X"81065156",
        X"56748938",
        X"83569439",
        X"81569039",
        X"7c51fa94",
        X"3f83c080",
        X"08881c0c",
        X"fd813975",
        X"83c0800c",
        X"903d0d04",
        X"f83d0d7a",
        X"7c595782",
        X"5483fe53",
        X"77527651",
        X"a3eb3f83",
        X"5683c080",
        X"0880ec38",
        X"81173377",
        X"3371882b",
        X"07565682",
        X"567482d4",
        X"d52e0981",
        X"0680d438",
        X"7554b653",
        X"77527651",
        X"a3bf3f83",
        X"c0800898",
        X"38811733",
        X"77337188",
        X"2b0783c0",
        X"80085256",
        X"56748182",
        X"c62eac38",
        X"825480d2",
        X"53775276",
        X"51a3963f",
        X"83c08008",
        X"98388117",
        X"33773371",
        X"882b0783",
        X"c0800852",
        X"56567481",
        X"82c62e83",
        X"38815675",
        X"83c0800c",
        X"8a3d0d04",
        X"eb3d0d67",
        X"5a800b83",
        X"c0900ca2",
        X"b83f83c0",
        X"80088106",
        X"55825674",
        X"83ef3874",
        X"75538f3d",
        X"70535759",
        X"feca3f83",
        X"c0800881",
        X"ff065776",
        X"812e0981",
        X"0680d438",
        X"905483be",
        X"53745275",
        X"51a2aa3f",
        X"83c08008",
        X"80c9388f",
        X"3d335574",
        X"802e80c9",
        X"3802bf05",
        X"33028405",
        X"be053371",
        X"982b7190",
        X"2b07028c",
        X"05bd0533",
        X"70882b72",
        X"07953d33",
        X"71077058",
        X"7b575e52",
        X"5e575957",
        X"fdee3f83",
        X"c0800881",
        X"ff065776",
        X"832e0981",
        X"06863881",
        X"5682f239",
        X"76802e86",
        X"38865682",
        X"e839a454",
        X"8d537852",
        X"7551a1c1",
        X"3f815683",
        X"c0800882",
        X"d43802be",
        X"05330284",
        X"05bd0533",
        X"71882b07",
        X"595d77ab",
        X"380280ce",
        X"05330284",
        X"0580cd05",
        X"3371982b",
        X"71902b07",
        X"973d3370",
        X"882b7207",
        X"02940580",
        X"cb053371",
        X"0754525e",
        X"57595602",
        X"b7053378",
        X"71290288",
        X"05b60533",
        X"028c05b5",
        X"05337188",
        X"2b07701d",
        X"707f8c05",
        X"0c5f5957",
        X"595d8e3d",
        X"33821b34",
        X"02b90533",
        X"903d3371",
        X"882b075a",
        X"5c78841b",
        X"2302bb05",
        X"33028405",
        X"ba053371",
        X"882b0756",
        X"5c74ab38",
        X"0280ca05",
        X"33028405",
        X"80c90533",
        X"71982b71",
        X"902b0796",
        X"3d337088",
        X"2b720702",
        X"940580c7",
        X"05337107",
        X"51525357",
        X"5e5c7476",
        X"31783179",
        X"842a903d",
        X"33547171",
        X"31535656",
        X"80d5a43f",
        X"83c08008",
        X"82057088",
        X"1c0c83c0",
        X"8008e08a",
        X"05565674",
        X"83dffe26",
        X"83388257",
        X"83fff676",
        X"27853883",
        X"57893986",
        X"5676802e",
        X"80db3876",
        X"7a347683",
        X"2e098106",
        X"b0380280",
        X"d6053302",
        X"840580d5",
        X"05337198",
        X"2b71902b",
        X"07993d33",
        X"70882b72",
        X"07029405",
        X"80d30533",
        X"71077f90",
        X"050c525e",
        X"57585686",
        X"39771b90",
        X"1b0c841a",
        X"228c1b08",
        X"1971842a",
        X"05941c0c",
        X"5d800b81",
        X"1b347983",
        X"c0900c80",
        X"567583c0",
        X"800c973d",
        X"0d04e93d",
        X"0d83c090",
        X"08568554",
        X"75802e81",
        X"8238800b",
        X"81173499",
        X"3de01146",
        X"6a548a3d",
        X"705458ec",
        X"0551f6e5",
        X"3f83c080",
        X"085483c0",
        X"800880df",
        X"38893d33",
        X"5473802e",
        X"913802ab",
        X"05337084",
        X"2a810651",
        X"5574802e",
        X"86388354",
        X"80c13976",
        X"51f4893f",
        X"83c08008",
        X"a0170c02",
        X"bf053302",
        X"8405be05",
        X"3371982b",
        X"71902b07",
        X"028c05bd",
        X"05337088",
        X"2b720795",
        X"3d337107",
        X"9c1c0c52",
        X"78981b0c",
        X"53565957",
        X"810b8117",
        X"34745473",
        X"83c0800c",
        X"993d0d04",
        X"f53d0d7d",
        X"7f617283",
        X"c090085a",
        X"5d5d595c",
        X"807b0c85",
        X"5775802e",
        X"81e03881",
        X"16338106",
        X"55845774",
        X"802e81d2",
        X"38913974",
        X"81173486",
        X"39800b81",
        X"17348157",
        X"81c0399c",
        X"16089817",
        X"08315574",
        X"78278338",
        X"74587780",
        X"2e81a938",
        X"98160870",
        X"83ff0656",
        X"577480cf",
        X"38821633",
        X"ff057789",
        X"2a067081",
        X"ff065a55",
        X"78a03876",
        X"8738a016",
        X"08558d39",
        X"a4160851",
        X"f0e93f83",
        X"c0800855",
        X"817527ff",
        X"a83874a4",
        X"170ca416",
        X"0851f283",
        X"3f83c080",
        X"085583c0",
        X"8008802e",
        X"ff893883",
        X"c0800819",
        X"a8170c98",
        X"160883ff",
        X"06848071",
        X"31515577",
        X"75278338",
        X"77557483",
        X"ffff0654",
        X"98160883",
        X"ff0653a8",
        X"16085279",
        X"577b8338",
        X"7b577651",
        X"9be73f83",
        X"c08008fe",
        X"d0389816",
        X"08159817",
        X"0c741a78",
        X"76317c08",
        X"177d0c59",
        X"5afed339",
        X"80577683",
        X"c0800c8d",
        X"3d0d04fa",
        X"3d0d7883",
        X"c0900855",
        X"56855573",
        X"802e81e3",
        X"38811433",
        X"81065384",
        X"5572802e",
        X"81d5389c",
        X"14085372",
        X"76278338",
        X"72569814",
        X"0857800b",
        X"98150c75",
        X"802e81b9",
        X"38821433",
        X"70892b56",
        X"5376802e",
        X"b7387452",
        X"ff165180",
        X"d0a53f83",
        X"c08008ff",
        X"18765470",
        X"53585380",
        X"d0953f83",
        X"c0800873",
        X"26963874",
        X"30707806",
        X"7098170c",
        X"777131a4",
        X"17085258",
        X"51538939",
        X"a0140870",
        X"a4160c53",
        X"747627b9",
        X"387251ee",
        X"d63f83c0",
        X"80085381",
        X"0b83c080",
        X"08278b38",
        X"88140883",
        X"c0800826",
        X"8838800b",
        X"811534b0",
        X"3983c080",
        X"08a4150c",
        X"98140815",
        X"98150c75",
        X"753156c4",
        X"39981408",
        X"16709816",
        X"0c735256",
        X"efc53f83",
        X"c080088c",
        X"3883c080",
        X"08811534",
        X"81559439",
        X"821433ff",
        X"0576892a",
        X"0683c080",
        X"0805a815",
        X"0c805574",
        X"83c0800c",
        X"883d0d04",
        X"ef3d0d63",
        X"56855583",
        X"c0900880",
        X"2e80d238",
        X"933df405",
        X"84170c64",
        X"53883d70",
        X"53765257",
        X"f1cf3f83",
        X"c0800855",
        X"83c08008",
        X"b438883d",
        X"33547380",
        X"2ea13802",
        X"a7053370",
        X"842a7081",
        X"06515555",
        X"83557380",
        X"2e973876",
        X"51eef53f",
        X"83c08008",
        X"88170c75",
        X"51efa63f",
        X"83c08008",
        X"557483c0",
        X"800c933d",
        X"0d04e43d",
        X"0d6ea13d",
        X"08405e85",
        X"5683c090",
        X"08802e84",
        X"85389e3d",
        X"f405841f",
        X"0c7e9838",
        X"7d51eef5",
        X"3f83c080",
        X"085683ee",
        X"39814181",
        X"f6398341",
        X"81f13993",
        X"3d7f9605",
        X"4159807f",
        X"8295055e",
        X"56756081",
        X"ff053483",
        X"41901e08",
        X"762e81d3",
        X"38a0547d",
        X"2270852b",
        X"83e00654",
        X"58901e08",
        X"52785197",
        X"f03f83c0",
        X"80084183",
        X"c08008ff",
        X"b8387833",
        X"5c7b802e",
        X"ffb4388b",
        X"193370bf",
        X"06718106",
        X"52435574",
        X"802e80de",
        X"387b81bf",
        X"0655748f",
        X"2480d338",
        X"9a193355",
        X"7480cb38",
        X"f31d7058",
        X"5d815675",
        X"8b2e0981",
        X"0685388e",
        X"568b3975",
        X"9a2e0981",
        X"0683389c",
        X"56781670",
        X"70810552",
        X"33713381",
        X"1a821a5f",
        X"5b525b55",
        X"74863879",
        X"77348539",
        X"80df7734",
        X"777b5757",
        X"7aa02e09",
        X"8106c038",
        X"81567b81",
        X"e5327030",
        X"709f2a51",
        X"51557bae",
        X"2e933874",
        X"802e8e38",
        X"61832a70",
        X"81065155",
        X"74802e97",
        X"387d51ed",
        X"df3f83c0",
        X"80084183",
        X"c0800887",
        X"38901e08",
        X"feaf3880",
        X"60347580",
        X"2e88387c",
        X"527f518f",
        X"963f6080",
        X"2e863880",
        X"0b901f0c",
        X"60566083",
        X"2e853860",
        X"81d03889",
        X"1f57901e",
        X"08802e81",
        X"a8388056",
        X"78167033",
        X"515574a0",
        X"2ea03874",
        X"852e0981",
        X"06843881",
        X"e5557477",
        X"70810559",
        X"34811670",
        X"81ff0657",
        X"55877627",
        X"d7388819",
        X"335574a0",
        X"2ea938ae",
        X"77708105",
        X"59348856",
        X"78167033",
        X"515574a0",
        X"2e953874",
        X"77708105",
        X"59348116",
        X"7081ff06",
        X"57558a76",
        X"27e2388b",
        X"19337f88",
        X"05349f19",
        X"339e1a33",
        X"71982b71",
        X"902b079d",
        X"1c337088",
        X"2b72079c",
        X"1e337107",
        X"640c5299",
        X"1d33981e",
        X"3371882b",
        X"07535153",
        X"57595674",
        X"7f840523",
        X"97193396",
        X"1a337188",
        X"2b075656",
        X"747f8605",
        X"23807734",
        X"7d51ebf0",
        X"3f83c080",
        X"08833270",
        X"30707207",
        X"9f2c83c0",
        X"80080652",
        X"5656961f",
        X"3355748a",
        X"38891f52",
        X"961f518d",
        X"a23f7583",
        X"c0800c9e",
        X"3d0d04f4",
        X"3d0d7e8f",
        X"3dec1156",
        X"56589053",
        X"f0155277",
        X"51e0d23f",
        X"83c08008",
        X"80d63878",
        X"902e0981",
        X"0680cd38",
        X"02ab0533",
        X"80fcb40b",
        X"80fcb433",
        X"5758568c",
        X"3974762e",
        X"8a388417",
        X"70335657",
        X"74f33876",
        X"33705755",
        X"74802eac",
        X"38821722",
        X"708a2b90",
        X"3dec0556",
        X"70555656",
        X"96800a52",
        X"7751e081",
        X"3f83c080",
        X"08863878",
        X"752e8538",
        X"80568539",
        X"81173356",
        X"7583c080",
        X"0c8e3d0d",
        X"04fc3d0d",
        X"76705255",
        X"8ca93f83",
        X"c0800815",
        X"ff055473",
        X"752e8e38",
        X"73335372",
        X"ae2e8638",
        X"ff1454ef",
        X"39775281",
        X"14518bc1",
        X"3f83c080",
        X"08307083",
        X"c0800807",
        X"802583c0",
        X"800c5386",
        X"3d0d04fc",
        X"3d0d7670",
        X"5255e6ee",
        X"3f83c080",
        X"08548153",
        X"83c08008",
        X"80c13874",
        X"51e6b13f",
        X"83c08008",
        X"80faa453",
        X"83c08008",
        X"5253ff91",
        X"3f83c080",
        X"08a13880",
        X"faa85272",
        X"51ff823f",
        X"83c08008",
        X"923880fa",
        X"ac527251",
        X"fef33f83",
        X"c0800880",
        X"2e833881",
        X"54735372",
        X"83c0800c",
        X"863d0d04",
        X"fc3d0d76",
        X"705255e6",
        X"8d3f83c0",
        X"80085481",
        X"5383c080",
        X"0880d138",
        X"7451e5d0",
        X"3f83c080",
        X"0880faa4",
        X"5383c080",
        X"085253fe",
        X"b03f83c0",
        X"8008b138",
        X"80faa852",
        X"7251fea1",
        X"3f83c080",
        X"08a23880",
        X"faac5272",
        X"51fe923f",
        X"83c08008",
        X"933883c3",
        X"9c085272",
        X"51fe823f",
        X"83c08008",
        X"802e8338",
        X"81547353",
        X"7283c080",
        X"0c863d0d",
        X"04fd3d0d",
        X"75705254",
        X"e59c3f81",
        X"5383c080",
        X"08983873",
        X"51e4e53f",
        X"83c38c08",
        X"5283c080",
        X"0851fdc9",
        X"3f83c080",
        X"08537283",
        X"c0800c85",
        X"3d0d04df",
        X"3d0da43d",
        X"0870525e",
        X"db833f83",
        X"c0800833",
        X"953d5654",
        X"73963880",
        X"ffd05274",
        X"5189b03f",
        X"9a397d52",
        X"7851de8b",
        X"3f84cc39",
        X"7d51dae9",
        X"3f83c080",
        X"08527451",
        X"da993f80",
        X"43804280",
        X"41804083",
        X"c3940852",
        X"943d7052",
        X"5de0f33f",
        X"83c08008",
        X"59800b83",
        X"c0800855",
        X"5b83c080",
        X"087b2e94",
        X"38811b74",
        X"525be3f5",
        X"3f83c080",
        X"085483c0",
        X"8008ee38",
        X"805aff5f",
        X"7909709f",
        X"2c7b065b",
        X"547a7a24",
        X"8438ff1b",
        X"5af61a70",
        X"09709f2c",
        X"72067bff",
        X"125a5a52",
        X"55558075",
        X"25953876",
        X"51e3ba3f",
        X"83c08008",
        X"76ff1858",
        X"55577380",
        X"24ed3874",
        X"7f2e8638",
        X"a2843f74",
        X"5f78ff1b",
        X"70585d58",
        X"807a2595",
        X"387751e3",
        X"903f83c0",
        X"800876ff",
        X"18585558",
        X"738024ed",
        X"38800b83",
        X"c7c40c80",
        X"0b83c7f0",
        X"0c80fab0",
        X"518daf3f",
        X"81800b83",
        X"c7f00c80",
        X"fab8518d",
        X"a13fa80b",
        X"83c7c40c",
        X"76802e80",
        X"e43883c7",
        X"c4087779",
        X"32703070",
        X"72078025",
        X"70872b83",
        X"c7f00c51",
        X"56785356",
        X"56e2c73f",
        X"83c08008",
        X"802e8838",
        X"80fac051",
        X"8ce83f76",
        X"51e2893f",
        X"83c08008",
        X"5280fb80",
        X"518cd73f",
        X"7651e291",
        X"3f83c080",
        X"0883c7c4",
        X"08555775",
        X"74258638",
        X"a81656f7",
        X"397583c7",
        X"c40c86f0",
        X"7624ff98",
        X"3887980b",
        X"83c7c40c",
        X"77802eb1",
        X"387751e1",
        X"c73f83c0",
        X"80087852",
        X"55e1e73f",
        X"80fac854",
        X"83c08008",
        X"8d388739",
        X"80763481",
        X"ec3980fa",
        X"80547453",
        X"735280fa",
        X"cc518bf6",
        X"3f805480",
        X"fad4518b",
        X"ed3f8114",
        X"5473a82e",
        X"098106ef",
        X"38868da0",
        X"519df73f",
        X"8052903d",
        X"70525880",
        X"c5993f83",
        X"52775180",
        X"c5913f62",
        X"81ab3861",
        X"802e8197",
        X"387b5473",
        X"ff2e9638",
        X"78802e81",
        X"86387851",
        X"e0eb3f83",
        X"c08008ff",
        X"155559e7",
        X"3978802e",
        X"80f13878",
        X"51e0e73f",
        X"83c08008",
        X"802efc8e",
        X"387851e0",
        X"af3f83c0",
        X"80085280",
        X"faa05184",
        X"833f83c0",
        X"8008bb38",
        X"7c5185bb",
        X"3f83c080",
        X"08ff0555",
        X"800b83c0",
        X"80082580",
        X"c838a33d",
        X"7505c405",
        X"70585676",
        X"33ff1858",
        X"5473af2e",
        X"fec23874",
        X"ff16ff18",
        X"58565473",
        X"8024e838",
        X"a4397851",
        X"dfd83f83",
        X"c0800852",
        X"7c5184db",
        X"3f933981",
        X"549f397f",
        X"10608829",
        X"057a0561",
        X"055afbf4",
        X"3962802e",
        X"fbb53880",
        X"52775180",
        X"c3d53f80",
        X"547383c0",
        X"800ca33d",
        X"0d04803d",
        X"0d9088b8",
        X"337081ff",
        X"0670842a",
        X"81327081",
        X"06515151",
        X"5170802e",
        X"8d38a80b",
        X"9088b834",
        X"b80b9088",
        X"b8347083",
        X"c0800c82",
        X"3d0d0480",
        X"3d0d9088",
        X"b8337081",
        X"ff067085",
        X"2a813270",
        X"81065151",
        X"51517080",
        X"2e8d3898",
        X"0b9088b8",
        X"34b80b90",
        X"88b83470",
        X"83c0800c",
        X"823d0d04",
        X"930b9088",
        X"bc34ff0b",
        X"9088a834",
        X"04ff3d0d",
        X"028f0533",
        X"52800b90",
        X"88bc348a",
        X"519b9b3f",
        X"df3f80f8",
        X"0b9088a0",
        X"34800b90",
        X"888834fa",
        X"12527190",
        X"88803480",
        X"0b908898",
        X"34719088",
        X"90349088",
        X"b8528072",
        X"34b87234",
        X"833d0d04",
        X"803d0d02",
        X"8b053351",
        X"709088b4",
        X"34febf3f",
        X"83c08008",
        X"802ef638",
        X"823d0d04",
        X"803d0d84",
        X"39a3e43f",
        X"fed93f83",
        X"c0800880",
        X"2ef33890",
        X"88b43370",
        X"81ff0683",
        X"c0800c51",
        X"823d0d04",
        X"803d0da3",
        X"0b9088bc",
        X"34ff0b90",
        X"88a83490",
        X"88b851a8",
        X"7134b871",
        X"34823d0d",
        X"04803d0d",
        X"9088bc33",
        X"70982b70",
        X"802583c0",
        X"800c5151",
        X"823d0d04",
        X"803d0d90",
        X"88b83370",
        X"81ff0670",
        X"832a8132",
        X"70810651",
        X"51515170",
        X"802ee838",
        X"b00b9088",
        X"b834b80b",
        X"9088b834",
        X"823d0d04",
        X"803d0d90",
        X"80ac0881",
        X"0683c080",
        X"0c823d0d",
        X"04fd3d0d",
        X"75775454",
        X"80732594",
        X"38737081",
        X"05553352",
        X"80fad851",
        X"87843fff",
        X"1353e939",
        X"853d0d04",
        X"fd3d0d75",
        X"77535473",
        X"33517089",
        X"38713351",
        X"70802ea1",
        X"38733372",
        X"33525372",
        X"71278538",
        X"ff519439",
        X"70732785",
        X"3881518b",
        X"39811481",
        X"135354d3",
        X"39805170",
        X"83c0800c",
        X"853d0d04",
        X"fd3d0d75",
        X"77545472",
        X"337081ff",
        X"06525270",
        X"802ea338",
        X"7181ff06",
        X"8114ffbf",
        X"12535452",
        X"70992689",
        X"38a01270",
        X"81ff0653",
        X"51717470",
        X"81055634",
        X"d2398074",
        X"34853d0d",
        X"04ffbd3d",
        X"0d80c63d",
        X"0852a53d",
        X"705254ff",
        X"b33f80c7",
        X"3d085285",
        X"3d705253",
        X"ffa63f72",
        X"527351fe",
        X"df3f80c5",
        X"3d0d04fe",
        X"3d0d7476",
        X"53537170",
        X"81055333",
        X"51707370",
        X"81055534",
        X"70f03884",
        X"3d0d04fe",
        X"3d0d7452",
        X"80723352",
        X"5370732e",
        X"8d388112",
        X"81147133",
        X"53545270",
        X"f5387283",
        X"c0800c84",
        X"3d0d04f6",
        X"3d0d7c7e",
        X"60625a5d",
        X"5b568059",
        X"81558539",
        X"747a2955",
        X"74527551",
        X"bbe93f83",
        X"c080087a",
        X"27ee3874",
        X"802e80dd",
        X"38745275",
        X"51bbd43f",
        X"83c08008",
        X"75537652",
        X"54bbd83f",
        X"83c08008",
        X"7a537552",
        X"56bbbc3f",
        X"83c08008",
        X"7930707b",
        X"079f2a70",
        X"77802407",
        X"51515455",
        X"72873883",
        X"c08008c5",
        X"38768118",
        X"b0165558",
        X"58897425",
        X"8b38b714",
        X"537a8538",
        X"80d71453",
        X"72783481",
        X"1959ff9f",
        X"39807734",
        X"8c3d0d04",
        X"f73d0d7b",
        X"7d7f6202",
        X"9005bb05",
        X"33575956",
        X"5a5ab058",
        X"728338a0",
        X"58757070",
        X"81055233",
        X"71595455",
        X"90398074",
        X"258e38ff",
        X"14777081",
        X"05593354",
        X"5472ef38",
        X"73ff1555",
        X"53807325",
        X"89387752",
        X"7951782d",
        X"ef397533",
        X"75575372",
        X"802e9038",
        X"72527951",
        X"782d7570",
        X"81055733",
        X"53ed398b",
        X"3d0d04ee",
        X"3d0d6466",
        X"69697070",
        X"81055233",
        X"5b4a5c5e",
        X"5e76802e",
        X"82f93876",
        X"a52e0981",
        X"0682e038",
        X"80704167",
        X"70708105",
        X"5233714a",
        X"59575f76",
        X"b02e0981",
        X"068c3875",
        X"70810557",
        X"33764857",
        X"815fd017",
        X"56758926",
        X"80da3876",
        X"675c5980",
        X"5c933977",
        X"8a2480c3",
        X"387b8a29",
        X"187b7081",
        X"055d335a",
        X"5cd01970",
        X"81ff0658",
        X"58897727",
        X"a438ff9f",
        X"197081ff",
        X"06ffa91b",
        X"5a515685",
        X"76279238",
        X"ffbf1970",
        X"81ff0651",
        X"56758526",
        X"8a38c919",
        X"58778025",
        X"ffb9387a",
        X"477b4078",
        X"81ff0657",
        X"7680e42e",
        X"80e53876",
        X"80e424a7",
        X"387680d8",
        X"2e818638",
        X"7680d824",
        X"90387680",
        X"2e81cc38",
        X"76a52e81",
        X"b63881b9",
        X"397680e3",
        X"2e818c38",
        X"81af3976",
        X"80f52e9b",
        X"387680f5",
        X"248b3876",
        X"80f32e81",
        X"81388199",
        X"397680f8",
        X"2e80ca38",
        X"818f3991",
        X"3d705557",
        X"80538a52",
        X"79841b71",
        X"08535b56",
        X"fc813f76",
        X"55ab3979",
        X"841b7108",
        X"943d705b",
        X"5b525b56",
        X"7580258c",
        X"38753056",
        X"ad783402",
        X"80c10557",
        X"76548053",
        X"8a527551",
        X"fbd53f77",
        X"557e54b8",
        X"39913d70",
        X"557780d8",
        X"32703070",
        X"80255651",
        X"58569052",
        X"79841b71",
        X"08535b57",
        X"fbb13f75",
        X"55db3979",
        X"841b8312",
        X"33545b56",
        X"98397984",
        X"1b710857",
        X"5b568054",
        X"7f537c52",
        X"7d51fc9c",
        X"3f873976",
        X"527d517c",
        X"2d667033",
        X"58810547",
        X"fd833994",
        X"3d0d0472",
        X"83c0940c",
        X"7183c098",
        X"0c04fb3d",
        X"0d883d70",
        X"70840552",
        X"08575475",
        X"5383c094",
        X"085283c0",
        X"980851fc",
        X"c63f873d",
        X"0d04ff3d",
        X"0d737008",
        X"53510293",
        X"05337234",
        X"70088105",
        X"710c833d",
        X"0d04fc3d",
        X"0d873d88",
        X"11557854",
        X"bed25351",
        X"fc993f80",
        X"52873d51",
        X"d13f863d",
        X"0d04fc3d",
        X"0d765574",
        X"83c3a008",
        X"2eaf3880",
        X"53745187",
        X"c63f83c0",
        X"800881ff",
        X"06ff1470",
        X"81ff0672",
        X"30709f2a",
        X"51525553",
        X"5472802e",
        X"843871dd",
        X"3873fe38",
        X"7483c3a0",
        X"0c863d0d",
        X"04ff3d0d",
        X"ff0b83c3",
        X"a00c84a5",
        X"3f815187",
        X"8a3f83c0",
        X"800881ff",
        X"065271ee",
        X"3881d33f",
        X"7183c080",
        X"0c833d0d",
        X"04fc3d0d",
        X"76028405",
        X"a2052202",
        X"8805a605",
        X"227a5455",
        X"5555ff82",
        X"3f72802e",
        X"a03883c3",
        X"b4143375",
        X"70810557",
        X"34811470",
        X"83ffff06",
        X"ff157083",
        X"ffff0656",
        X"525552dd",
        X"39800b83",
        X"c0800c86",
        X"3d0d04fc",
        X"3d0d7678",
        X"7a115653",
        X"55805371",
        X"742e9338",
        X"74135170",
        X"3383c3b4",
        X"13348112",
        X"81145452",
        X"ea39800b",
        X"83c0800c",
        X"863d0d04",
        X"fd3d0d90",
        X"5483c3a0",
        X"085186f9",
        X"3f83c080",
        X"0881ff06",
        X"ff157130",
        X"71307073",
        X"079f2a72",
        X"9f2a0652",
        X"55525553",
        X"72db3885",
        X"3d0d0480",
        X"3d0d83c3",
        X"ac081083",
        X"c3a40807",
        X"9080a80c",
        X"823d0d04",
        X"800b83c3",
        X"ac0ce43f",
        X"04810b83",
        X"c3ac0cdb",
        X"3f04ed3f",
        X"047183c3",
        X"a80c0480",
        X"3d0d8051",
        X"f43f810b",
        X"83c3ac0c",
        X"810b83c3",
        X"a40cffbb",
        X"3f823d0d",
        X"04803d0d",
        X"72307074",
        X"07802583",
        X"c3a40c51",
        X"ffa53f82",
        X"3d0d0480",
        X"3d0d028b",
        X"05339080",
        X"a40c9080",
        X"a8087081",
        X"06515170",
        X"f5389080",
        X"a4087081",
        X"ff0683c0",
        X"800c5182",
        X"3d0d0480",
        X"3d0d81ff",
        X"51d13f83",
        X"c0800881",
        X"ff0683c0",
        X"800c823d",
        X"0d04803d",
        X"0d73902b",
        X"73079080",
        X"b40c823d",
        X"0d0404fb",
        X"3d0d7802",
        X"84059f05",
        X"3370982b",
        X"55575572",
        X"80259b38",
        X"7580ff06",
        X"56805280",
        X"f751e03f",
        X"83c08008",
        X"81ff0654",
        X"73812680",
        X"ff388051",
        X"fee73fff",
        X"a23f8151",
        X"fedf3fff",
        X"9a3f7551",
        X"feed3f74",
        X"982a51fe",
        X"e63f7490",
        X"2a7081ff",
        X"065253fe",
        X"da3f7488",
        X"2a7081ff",
        X"065253fe",
        X"ce3f7481",
        X"ff0651fe",
        X"c63f8155",
        X"7580c02e",
        X"09810686",
        X"38819555",
        X"8d397580",
        X"c82e0981",
        X"06843881",
        X"87557451",
        X"fea53f8a",
        X"55fec83f",
        X"83c08008",
        X"81ff0670",
        X"982b5454",
        X"7280258c",
        X"38ff1570",
        X"81ff0656",
        X"5374e238",
        X"7383c080",
        X"0c873d0d",
        X"04fa3d0d",
        X"fdc53f80",
        X"51fdda3f",
        X"8a54fe93",
        X"3fff1470",
        X"81ff0655",
        X"5373f338",
        X"73745355",
        X"80c051fe",
        X"a63f83c0",
        X"800881ff",
        X"06547381",
        X"2e098106",
        X"82a43883",
        X"aa5280c8",
        X"51fe8c3f",
        X"83c08008",
        X"81ff0653",
        X"72812e09",
        X"810681ad",
        X"38745488",
        X"3d7405fc",
        X"0553fdc7",
        X"3f83c080",
        X"08733481",
        X"147081ff",
        X"06555383",
        X"7427e438",
        X"029a0533",
        X"5372812e",
        X"09810681",
        X"dd38029b",
        X"05335380",
        X"ce905472",
        X"81aa2e8d",
        X"3881cb39",
        X"80e4518b",
        X"c53fff14",
        X"5473802e",
        X"81bc3882",
        X"0a5281e9",
        X"51fda43f",
        X"83c08008",
        X"81ff0653",
        X"72de3872",
        X"5280fa51",
        X"fd913f83",
        X"c0800881",
        X"ff065372",
        X"81943872",
        X"54883d74",
        X"05fc0553",
        X"fcd13f83",
        X"c0800873",
        X"34811470",
        X"81ff0655",
        X"53837427",
        X"e438873d",
        X"3370862a",
        X"70810651",
        X"54568c55",
        X"7280e338",
        X"845580de",
        X"39745281",
        X"e951fcc7",
        X"3f83c080",
        X"0881ff06",
        X"53825581",
        X"e9568173",
        X"27863873",
        X"5580c156",
        X"80ce9054",
        X"8a3980e4",
        X"518ab33f",
        X"ff145473",
        X"802ea938",
        X"80527551",
        X"fc953f83",
        X"c0800881",
        X"ff065372",
        X"e1388480",
        X"5280d051",
        X"fc813f83",
        X"c0800881",
        X"ff065372",
        X"802e8338",
        X"80557483",
        X"c3b03480",
        X"51fb823f",
        X"fbbd3f88",
        X"3d0d04fb",
        X"3d0d7754",
        X"800b83c3",
        X"b0337083",
        X"2a708106",
        X"51555755",
        X"72752e09",
        X"81068538",
        X"73892b54",
        X"735280d1",
        X"51fbb83f",
        X"83c08008",
        X"81ff0653",
        X"72bd3882",
        X"b8c054fa",
        X"fe3f83c0",
        X"800881ff",
        X"06537281",
        X"ff2e0981",
        X"068938ff",
        X"145473e7",
        X"389f3972",
        X"81fe2e09",
        X"81069638",
        X"83c7b452",
        X"83c3b451",
        X"fae83ffa",
        X"ce3ffacb",
        X"3f833981",
        X"558051fa",
        X"843ffabf",
        X"3f7481ff",
        X"0683c080",
        X"0c873d0d",
        X"04fb3d0d",
        X"7783c3b4",
        X"56548151",
        X"f9e73f83",
        X"c3b03370",
        X"832a7081",
        X"06515456",
        X"72853873",
        X"892b5473",
        X"5280d851",
        X"fab13f83",
        X"c0800881",
        X"ff065372",
        X"80e43881",
        X"ff51f9cf",
        X"3f81fe51",
        X"f9c93f84",
        X"80537470",
        X"81055633",
        X"51f9bc3f",
        X"ff137083",
        X"ffff0651",
        X"5372eb38",
        X"7251f9ab",
        X"3f7251f9",
        X"a63ff9cb",
        X"3f83c080",
        X"089f0653",
        X"a7885472",
        X"852e8c38",
        X"993980e4",
        X"5187eb3f",
        X"ff1454f9",
        X"ae3f83c0",
        X"800881ff",
        X"2e843873",
        X"e9388051",
        X"f8df3ff9",
        X"9a3f800b",
        X"83c0800c",
        X"873d0d04",
        X"7183c7b8",
        X"0c888080",
        X"0b83c7b4",
        X"0c848080",
        X"0b83c7bc",
        X"0c04fd3d",
        X"0d777017",
        X"557705ff",
        X"1a535371",
        X"ff2e9438",
        X"73708105",
        X"55335170",
        X"73708105",
        X"5534ff12",
        X"52e93985",
        X"3d0d04fb",
        X"3d0d87a6",
        X"810b83c7",
        X"b8085656",
        X"753383a6",
        X"801634a0",
        X"5483a080",
        X"5383c7b8",
        X"085283c7",
        X"b40851ff",
        X"b13fa054",
        X"83a48053",
        X"83c7b808",
        X"5283c7b4",
        X"0851ff9e",
        X"3f905483",
        X"a8805383",
        X"c7b80852",
        X"83c7b408",
        X"51ff8b3f",
        X"a0538052",
        X"83c7bc08",
        X"83a08005",
        X"5186bc3f",
        X"a0538052",
        X"83c7bc08",
        X"83a48005",
        X"5186ac3f",
        X"90538052",
        X"83c7bc08",
        X"83a88005",
        X"51869c3f",
        X"ff763483",
        X"a0805480",
        X"5383c7b8",
        X"085283c7",
        X"bc0851fe",
        X"c53f80d0",
        X"805483b0",
        X"805383c7",
        X"b8085283",
        X"c7bc0851",
        X"feb03f87",
        X"e13fa254",
        X"805383c7",
        X"bc088c80",
        X"055280fd",
        X"a851fe9a",
        X"3f860b87",
        X"a8833480",
        X"0b87a882",
        X"34800b87",
        X"a09a34af",
        X"0b87a096",
        X"34bf0b87",
        X"a0973480",
        X"0b87a098",
        X"349f0b87",
        X"a0993480",
        X"0b87a09b",
        X"34e00b87",
        X"a88934a2",
        X"0b87a880",
        X"34830b87",
        X"a48f3482",
        X"0b87a881",
        X"34873d0d",
        X"04fc3d0d",
        X"83a08054",
        X"805383c7",
        X"bc085283",
        X"c7b80851",
        X"fdb83f80",
        X"d0805483",
        X"b0805383",
        X"c7bc0852",
        X"83c7b808",
        X"51fda33f",
        X"a05483a0",
        X"805383c7",
        X"bc085283",
        X"c7b80851",
        X"fd903fa0",
        X"5483a480",
        X"5383c7bc",
        X"085283c7",
        X"b80851fc",
        X"fd3f9054",
        X"83a88053",
        X"83c7bc08",
        X"5283c7b8",
        X"0851fcea",
        X"3f83c7b8",
        X"085583a6",
        X"80153387",
        X"a6813486",
        X"3d0d04fa",
        X"3d0d7870",
        X"5255c0ca",
        X"3f83ffff",
        X"0b83c080",
        X"0825a938",
        X"7451c0cb",
        X"3f83c080",
        X"089e3883",
        X"c0800857",
        X"883dfc05",
        X"54848080",
        X"5383c7b8",
        X"08527451",
        X"ffbdfd3f",
        X"ffbdc33f",
        X"883d0d04",
        X"fa3d0d78",
        X"705255c0",
        X"893f83ff",
        X"ff0b83c0",
        X"80082597",
        X"38805788",
        X"3dfc0554",
        X"84808053",
        X"83c7b808",
        X"527451ff",
        X"befb3f88",
        X"3d0d0480",
        X"3d0d9080",
        X"90088106",
        X"83c0800c",
        X"823d0d04",
        X"ff3d0d90",
        X"80907008",
        X"70fe0676",
        X"07720c52",
        X"52833d0d",
        X"04803d0d",
        X"90809008",
        X"70812c81",
        X"0683c080",
        X"0c51823d",
        X"0d04ff3d",
        X"0d908090",
        X"700870fd",
        X"06761007",
        X"720c5252",
        X"833d0d04",
        X"803d0d90",
        X"80900870",
        X"822cbf06",
        X"83c0800c",
        X"51823d0d",
        X"04ff3d0d",
        X"90809070",
        X"0870fe83",
        X"0676822b",
        X"07720c52",
        X"52833d0d",
        X"04803d0d",
        X"90809008",
        X"70882c87",
        X"0683c080",
        X"0c51823d",
        X"0d04ff3d",
        X"0d908090",
        X"700870f1",
        X"ff067688",
        X"2b07720c",
        X"5252833d",
        X"0d04803d",
        X"0d908090",
        X"0870912c",
        X"bf0683c0",
        X"800c5182",
        X"3d0d04ff",
        X"3d0d9080",
        X"90700870",
        X"fc87ffff",
        X"0676912b",
        X"07720c52",
        X"52833d0d",
        X"04803d0d",
        X"90809008",
        X"70992c81",
        X"0683c080",
        X"0c51823d",
        X"0d04ff3d",
        X"0d908090",
        X"700870ff",
        X"bf0a0676",
        X"992b0772",
        X"0c525283",
        X"3d0d0480",
        X"3d0d9080",
        X"80087088",
        X"2c810683",
        X"c0800c51",
        X"823d0d04",
        X"803d0d90",
        X"80800870",
        X"892c8106",
        X"83c0800c",
        X"51823d0d",
        X"04803d0d",
        X"90808008",
        X"708a2c81",
        X"0683c080",
        X"0c51823d",
        X"0d04803d",
        X"0d908080",
        X"08708b2c",
        X"810683c0",
        X"800c5182",
        X"3d0d0480",
        X"3d0d9080",
        X"80087092",
        X"2c810683",
        X"c0800c51",
        X"823d0d04",
        X"803d0d90",
        X"80800870",
        X"8c2cbf06",
        X"83c0800c",
        X"51823d0d",
        X"04803d0d",
        X"90808408",
        X"870683c0",
        X"800c823d",
        X"0d04fe3d",
        X"0d7481e6",
        X"29872a90",
        X"80a00c84",
        X"3d0d04fe",
        X"3d0d7575",
        X"ff195353",
        X"5370ff2e",
        X"8d387272",
        X"70810554",
        X"34ff1151",
        X"f039843d",
        X"0d04fe3d",
        X"0d7575ff",
        X"19535353",
        X"70ff2e8d",
        X"38727270",
        X"8405540c",
        X"ff1151f0",
        X"39843d0d",
        X"04fe3d0d",
        X"84808053",
        X"80528880",
        X"0a51ffb3",
        X"3f818080",
        X"53805282",
        X"800a51c6",
        X"3f843d0d",
        X"04803d0d",
        X"8151fc84",
        X"3f72802e",
        X"90388051",
        X"fdd83fcd",
        X"3f83c7c0",
        X"3351fdce",
        X"3f8151fc",
        X"953f8051",
        X"fc903f80",
        X"51fbe13f",
        X"823d0d04",
        X"fd3d0d75",
        X"52805480",
        X"ff722588",
        X"38810bff",
        X"80135354",
        X"ffbf1251",
        X"70992686",
        X"38e01252",
        X"b039ff9f",
        X"12519971",
        X"27a738d0",
        X"12e01354",
        X"51708926",
        X"85387252",
        X"9839728f",
        X"26853872",
        X"528f3971",
        X"ba2e0981",
        X"0685389a",
        X"52833980",
        X"5273802e",
        X"85388180",
        X"12527181",
        X"ff0683c0",
        X"800c853d",
        X"0d04803d",
        X"0d84d8c0",
        X"51807170",
        X"81055334",
        X"7084e0c0",
        X"2e098106",
        X"f038823d",
        X"0d04fe3d",
        X"0d029705",
        X"3351fef4",
        X"3f83c080",
        X"0881ff06",
        X"83c7c408",
        X"54528073",
        X"249b3883",
        X"c7ec0813",
        X"7283c7f0",
        X"08075353",
        X"71733483",
        X"c7c40881",
        X"0583c7c4",
        X"0c843d0d",
        X"04fa3d0d",
        X"82800a1b",
        X"55805788",
        X"3dfc0554",
        X"79537452",
        X"7851ffb8",
        X"ec3f883d",
        X"0d04fe3d",
        X"0d83c7dc",
        X"08527451",
        X"ffbfcf3f",
        X"83c08008",
        X"8c387653",
        X"755283c7",
        X"dc0851c5",
        X"3f843d0d",
        X"04fe3d0d",
        X"83c7dc08",
        X"53755274",
        X"51ffba8d",
        X"3f83c080",
        X"088d3877",
        X"53765283",
        X"c7dc0851",
        X"ff9f3f84",
        X"3d0d04fe",
        X"3d0d83c7",
        X"dc0851ff",
        X"b9803f83",
        X"c0800881",
        X"80802e09",
        X"81068838",
        X"83c18080",
        X"539c3983",
        X"c7dc0851",
        X"ffb8e33f",
        X"83c08008",
        X"80d0802e",
        X"09810693",
        X"3883c1b0",
        X"805383c0",
        X"80085283",
        X"c7dc0851",
        X"fed33f84",
        X"3d0d04ed",
        X"3d0d8044",
        X"80438042",
        X"80418070",
        X"5a5bfde6",
        X"3f800b83",
        X"c7c40c80",
        X"0b83c7f0",
        X"0c80fae0",
        X"51e9b33f",
        X"81800b83",
        X"c7f00c80",
        X"fae451e9",
        X"a53f81c8",
        X"0b83c7c4",
        X"0c783070",
        X"7a078025",
        X"70872b83",
        X"c7f00c51",
        X"5583c7dc",
        X"0851ffb4",
        X"f03f83c0",
        X"80085280",
        X"faec51e8",
        X"f93f8298",
        X"0b83c7c4",
        X"0c810b83",
        X"c7c85b58",
        X"83c7c408",
        X"79793270",
        X"30707207",
        X"80257087",
        X"2b83c7f0",
        X"0c51578e",
        X"3d7055ff",
        X"1b545757",
        X"5791d13f",
        X"79708405",
        X"5b0851ff",
        X"b4a73f74",
        X"5483c080",
        X"08537752",
        X"80faf451",
        X"e8ac3fa8",
        X"1783c7c4",
        X"0c811858",
        X"77852e09",
        X"8106ffb0",
        X"3883b80b",
        X"83c7c40c",
        X"78853270",
        X"30707207",
        X"80257087",
        X"2b83c7f0",
        X"0c515656",
        X"f8ac3f80",
        X"fb845583",
        X"c0800880",
        X"2e8f3883",
        X"c7d80851",
        X"ffb3d23f",
        X"83c08008",
        X"55745280",
        X"fb8c51e7",
        X"d93f8580",
        X"0b83c7c4",
        X"0c788632",
        X"70307072",
        X"07802570",
        X"872b83c7",
        X"f00c5156",
        X"80fb9852",
        X"56e7b73f",
        X"868da051",
        X"f9cc3ff8",
        X"f93f83c0",
        X"8008f838",
        X"83c08008",
        X"52913d70",
        X"5255a0e3",
        X"3f835274",
        X"51a0dc3f",
        X"63557482",
        X"97386119",
        X"59788025",
        X"85388659",
        X"90398679",
        X"25853874",
        X"59873978",
        X"862681f6",
        X"3878822b",
        X"5580fa84",
        X"15080460",
        X"87386280",
        X"2e81e338",
        X"83c39008",
        X"83c38c0c",
        X"aedd0b83",
        X"c3940c83",
        X"c7dc0851",
        X"d7a53ffc",
        X"a23f81c6",
        X"39605680",
        X"76259838",
        X"ad8b0b83",
        X"c3940c83",
        X"c7c41570",
        X"085255d7",
        X"863f7408",
        X"52923975",
        X"80259238",
        X"83c7c415",
        X"0851ffb2",
        X"923f8052",
        X"ff1951b8",
        X"3962802e",
        X"818c3883",
        X"c7c41570",
        X"0883c7c8",
        X"08720c83",
        X"c7c80cff",
        X"1a705351",
        X"558db53f",
        X"83c08008",
        X"5680518d",
        X"ab3f83c0",
        X"80085274",
        X"5189c43f",
        X"75528051",
        X"89bd3f80",
        X"d5396055",
        X"807525b6",
        X"3883c39c",
        X"0883c38c",
        X"0caedd0b",
        X"83c3940c",
        X"83c7d808",
        X"51d6903f",
        X"83c7d808",
        X"51d2c03f",
        X"83c08008",
        X"81ff0670",
        X"5255f5e3",
        X"3f74802e",
        X"9d388155",
        X"a1397480",
        X"25943883",
        X"c7d80851",
        X"ffb1843f",
        X"8051f5c7",
        X"3f843962",
        X"87387a80",
        X"2efbaf38",
        X"80557483",
        X"c0800c95",
        X"3d0d04fe",
        X"3d0d7476",
        X"ff195353",
        X"5370ff2e",
        X"92387170",
        X"81055333",
        X"73708105",
        X"5534ff11",
        X"51eb3984",
        X"3d0d04f5",
        X"3d0df5cf",
        X"3f83c080",
        X"08802e86",
        X"38805182",
        X"dd39f5d4",
        X"3f83c080",
        X"0882d138",
        X"f5f43f83",
        X"c0800880",
        X"2e819738",
        X"805c805b",
        X"805a8059",
        X"8151f3a8",
        X"3f8051f5",
        X"813fef9f",
        X"3f800b83",
        X"c7c40cfa",
        X"aa3f83c0",
        X"80085480",
        X"528d3df0",
        X"05519dbb",
        X"3ff5bb3f",
        X"83c08008",
        X"f838ff0b",
        X"83c7c40c",
        X"f0ff3f73",
        X"82823883",
        X"c7c03351",
        X"f4c83f73",
        X"51f2e53f",
        X"82cd3983",
        X"c7c80851",
        X"ffafc03f",
        X"80528051",
        X"87a53f83",
        X"c7cc0851",
        X"ffafb03f",
        X"80528151",
        X"87953f80",
        X"c45383c7",
        X"e8085283",
        X"c7d80851",
        X"feb13f83",
        X"c7d80851",
        X"d0a93f83",
        X"c0800851",
        X"f3d13f81",
        X"8e39f4bd",
        X"3f83c080",
        X"08802e81",
        X"ab388151",
        X"f28e3f80",
        X"51f3e73f",
        X"ee853fad",
        X"ec0b83c3",
        X"940c83c7",
        X"e80851d3",
        X"be3f83c0",
        X"80085883",
        X"c0800880",
        X"2e80d838",
        X"f4b13f83",
        X"c0800883",
        X"c39c0853",
        X"83c7e808",
        X"5257d0d5",
        X"3f83c080",
        X"08feec38",
        X"76567680",
        X"2e833881",
        X"5683c7d8",
        X"0851ffae",
        X"a23f8051",
        X"f2e53f75",
        X"842983c7",
        X"c8057008",
        X"555580c4",
        X"5383c7e8",
        X"08527351",
        X"fd9d3f74",
        X"08527551",
        X"85e93f76",
        X"ff9438f3",
        X"c53f83c0",
        X"8008f838",
        X"f3d13f83",
        X"c08008f8",
        X"38ff0b83",
        X"c7c40cef",
        X"803f7780",
        X"2e80dc38",
        X"8151f4e1",
        X"3f80d439",
        X"f3b13f83",
        X"c0800880",
        X"2e80c838",
        X"f3ba3f83",
        X"c0800890",
        X"2e098106",
        X"ba3883c7",
        X"c80883c7",
        X"cc0883c7",
        X"c80c83c7",
        X"cc0c8051",
        X"88ea3f83",
        X"c0800854",
        X"815188e0",
        X"3f83c080",
        X"08528051",
        X"84f93f73",
        X"52815184",
        X"f23ff2e7",
        X"3f83c080",
        X"08f83880",
        X"54f2dc3f",
        X"83c08008",
        X"742e8338",
        X"81547351",
        X"f0823f8d",
        X"3d0d04fb",
        X"3d0d800b",
        X"83c7c034",
        X"90808052",
        X"86848080",
        X"51ffb0e3",
        X"3f83c080",
        X"0881ae38",
        X"88a43f80",
        X"ffc051ff",
        X"b5a23f83",
        X"c0800855",
        X"9c800a54",
        X"80c08053",
        X"80fba052",
        X"83c08008",
        X"51f5de3f",
        X"83c7dc08",
        X"5380fbb0",
        X"527451ff",
        X"afeb3f83",
        X"c0800880",
        X"2e963883",
        X"c7dc0853",
        X"80fbbc52",
        X"7451ffaf",
        X"d43f83c0",
        X"80088438",
        X"f5d53f83",
        X"c7e00853",
        X"80fbcc52",
        X"7451ffaf",
        X"bc3f83c0",
        X"8008b638",
        X"873dfc05",
        X"54848080",
        X"5386a880",
        X"805283c7",
        X"e00851ff",
        X"adc73f83",
        X"c0800893",
        X"38758480",
        X"802e0981",
        X"06893881",
        X"0b83c7c0",
        X"34873980",
        X"0b83c7c0",
        X"3483c7c0",
        X"3351f09a",
        X"3f8151f2",
        X"ac3f9599",
        X"3f8151f2",
        X"a43f8151",
        X"facd3ffa",
        X"3983c08c",
        X"080283c0",
        X"8c0cfb3d",
        X"0d0280fb",
        X"d80b83c3",
        X"900c80fb",
        X"dc0b83c3",
        X"880c80fb",
        X"e00b83c3",
        X"9c0c80fb",
        X"e40b83c3",
        X"980c83c0",
        X"8c08fc05",
        X"0c800b83",
        X"c7c80b83",
        X"c08c08f8",
        X"050c83c0",
        X"8c08f405",
        X"0cffadcf",
        X"3f83c080",
        X"088605fc",
        X"0683c08c",
        X"08f0050c",
        X"0283c08c",
        X"08f00508",
        X"310d833d",
        X"7083c08c",
        X"08f80508",
        X"70840583",
        X"c08c08f8",
        X"050c0c51",
        X"ffaa903f",
        X"83c08c08",
        X"f4050881",
        X"0583c08c",
        X"08f4050c",
        X"83c08c08",
        X"f4050889",
        X"2e098106",
        X"ffab3886",
        X"94808051",
        X"e8c23fff",
        X"0b83c7c4",
        X"0c800b83",
        X"c7f00c84",
        X"d8c00b83",
        X"c7ec0c81",
        X"51ece93f",
        X"8151ed8e",
        X"3f8051ed",
        X"893fed9c",
        X"3f83c080",
        X"088b3881",
        X"51eda63f",
        X"8251edce",
        X"3f8051ed",
        X"f63f8051",
        X"eea03f80",
        X"d2ee5280",
        X"51dd983f",
        X"fcb93f83",
        X"c08c08fc",
        X"05080d80",
        X"0b83c080",
        X"0c873d0d",
        X"83c08c0c",
        X"04803d0d",
        X"81ff5180",
        X"0b83c7fc",
        X"1234ff11",
        X"5170f438",
        X"823d0d04",
        X"ff3d0d73",
        X"70335351",
        X"81113371",
        X"34718112",
        X"34833d0d",
        X"04fb3d0d",
        X"77795656",
        X"80707155",
        X"55527175",
        X"25ac3875",
        X"13703370",
        X"147081ff",
        X"06555151",
        X"51717427",
        X"89388112",
        X"7081ff06",
        X"53517181",
        X"147083ff",
        X"ff065552",
        X"54747324",
        X"d6387183",
        X"c0800c87",
        X"3d0d04f4",
        X"3d0d7e60",
        X"5955805d",
        X"8075822b",
        X"7183ca9c",
        X"120c83ca",
        X"b0175b5b",
        X"57767934",
        X"77772e83",
        X"b7387652",
        X"7751ffaa",
        X"9c3f8e3d",
        X"fc055490",
        X"5383ca84",
        X"527751ff",
        X"a9d73f7c",
        X"5675902e",
        X"09810683",
        X"933883ca",
        X"8451fed8",
        X"3f83ca86",
        X"51fed13f",
        X"83ca8851",
        X"feca3f76",
        X"83ca940c",
        X"7751ffa7",
        X"9c3f80fa",
        X"a85283c0",
        X"800851c9",
        X"bc3f83c0",
        X"8008812e",
        X"09810680",
        X"d4387683",
        X"caac0c82",
        X"0b83ca84",
        X"34ff960b",
        X"83ca8534",
        X"7751ffa9",
        X"e93f83c0",
        X"80085583",
        X"c0800877",
        X"25883883",
        X"c080088f",
        X"05557484",
        X"2c7083ff",
        X"ff067088",
        X"2a585155",
        X"7583ca86",
        X"347483ca",
        X"87347683",
        X"ca8834ff",
        X"800b83ca",
        X"89348190",
        X"3983ca84",
        X"3383ca85",
        X"3371882b",
        X"07565b74",
        X"83ffff2e",
        X"09810680",
        X"e838fe80",
        X"0b83caac",
        X"0c810b83",
        X"ca940cff",
        X"0b83ca84",
        X"34ff0b83",
        X"ca853477",
        X"51ffa8f6",
        X"3f83c080",
        X"0883cab4",
        X"0c83c080",
        X"085583c0",
        X"80088025",
        X"883883c0",
        X"80088f05",
        X"5574842c",
        X"7083ffff",
        X"0670882a",
        X"58515575",
        X"83ca8634",
        X"7483ca87",
        X"347683ca",
        X"8834ff80",
        X"0b83ca89",
        X"34810b83",
        X"ca9334a5",
        X"39748596",
        X"2e098106",
        X"80fe3875",
        X"83caac0c",
        X"7751ffa8",
        X"aa3f83ca",
        X"933383c0",
        X"80080755",
        X"7483ca93",
        X"3483ca93",
        X"33810655",
        X"74802e83",
        X"38845783",
        X"ca883383",
        X"ca893371",
        X"882b0756",
        X"5c748180",
        X"2e098106",
        X"a13883ca",
        X"863383ca",
        X"87337188",
        X"2b07565b",
        X"ad807527",
        X"87387682",
        X"07579c39",
        X"76810757",
        X"96397482",
        X"802e0981",
        X"06873876",
        X"83075787",
        X"397481ff",
        X"268a3877",
        X"83ca9c1b",
        X"0c767934",
        X"8e3d0d04",
        X"803d0d72",
        X"842983ca",
        X"9c057008",
        X"83c0800c",
        X"51823d0d",
        X"0404fe3d",
        X"0d83c09c",
        X"08873881",
        X"0b83c09c",
        X"0c800b83",
        X"ca800c80",
        X"0b83c9fc",
        X"0cff0b83",
        X"c7f80ca8",
        X"0b83ca98",
        X"0cae51ce",
        X"e83f800b",
        X"83ca9c54",
        X"52807370",
        X"8405550c",
        X"81125271",
        X"842e0981",
        X"06ef3884",
        X"3d0d04fe",
        X"3d0d7402",
        X"84059605",
        X"22535371",
        X"802e9638",
        X"72708105",
        X"543351ce",
        X"f33fff12",
        X"7083ffff",
        X"065152e7",
        X"39843d0d",
        X"04fe3d0d",
        X"02920522",
        X"5382ac51",
        X"e9c03f80",
        X"c351ced0",
        X"3f819651",
        X"e9b43f72",
        X"5283c7fc",
        X"51ffb43f",
        X"725283c7",
        X"fc51faa9",
        X"3f83c080",
        X"0881ff06",
        X"51cead3f",
        X"843d0d04",
        X"fc3d0d76",
        X"78718429",
        X"83ca9c05",
        X"70085153",
        X"5353709e",
        X"3880ce72",
        X"3480cf0b",
        X"81133480",
        X"ce0b8213",
        X"3480c50b",
        X"83133470",
        X"84133480",
        X"e73983ca",
        X"b0133354",
        X"80d27234",
        X"73822a70",
        X"81065151",
        X"80cf5370",
        X"843880d7",
        X"53728113",
        X"34a00b82",
        X"13347383",
        X"06517081",
        X"2e9e3870",
        X"81248838",
        X"70802e8f",
        X"389f3970",
        X"822e9238",
        X"70832e92",
        X"38933980",
        X"d8558e39",
        X"80d35589",
        X"3980cd55",
        X"843980c4",
        X"55748313",
        X"3480c40b",
        X"84133480",
        X"0b851334",
        X"863d0d04",
        X"803d0de7",
        X"e03f83c0",
        X"80088429",
        X"80ff8005",
        X"700883c0",
        X"800c5182",
        X"3d0d04ff",
        X"3d0d83ca",
        X"9808a82e",
        X"0981068d",
        X"38d63f83",
        X"c0800883",
        X"ca980c87",
        X"39a80b83",
        X"ca980c83",
        X"ca980886",
        X"057081ff",
        X"065252cc",
        X"803f833d",
        X"0d04fb3d",
        X"0d775689",
        X"39f0bc3f",
        X"8351e79a",
        X"3fcdcd3f",
        X"83c08008",
        X"802eee38",
        X"83ca9808",
        X"86057081",
        X"ff065253",
        X"cbd33f81",
        X"0b9088d4",
        X"34f0943f",
        X"8351e6f2",
        X"3f9088d4",
        X"337081ff",
        X"06555373",
        X"802eea38",
        X"73862a70",
        X"81065153",
        X"72ffbe38",
        X"73982b53",
        X"80732480",
        X"de38ccbd",
        X"3f83c080",
        X"085583c0",
        X"800880cf",
        X"38751575",
        X"822b5454",
        X"9088c013",
        X"33743481",
        X"15557485",
        X"2e098106",
        X"e8387533",
        X"83c7fc34",
        X"81163383",
        X"c7fd3482",
        X"163383c7",
        X"fe348316",
        X"3383c7ff",
        X"34845283",
        X"c7fc51f7",
        X"883f83c0",
        X"800881ff",
        X"06841733",
        X"55537274",
        X"2e8738fe",
        X"923ffed1",
        X"3980e451",
        X"e5e43f87",
        X"3d0d04ff",
        X"b23d0d80",
        X"d03df805",
        X"51feab3f",
        X"83ca8008",
        X"810583ca",
        X"800c80ce",
        X"3d33cf11",
        X"7081ff06",
        X"51565674",
        X"83268986",
        X"38758f06",
        X"ff055675",
        X"83c7f808",
        X"2e9b3875",
        X"83269638",
        X"7583c7f8",
        X"0c758429",
        X"83ca9c05",
        X"70085355",
        X"7551f6db",
        X"3f807624",
        X"88e23875",
        X"842983ca",
        X"9c055574",
        X"08802e88",
        X"d33883c7",
        X"f8088429",
        X"83ca9c05",
        X"70080288",
        X"0582b505",
        X"33525a55",
        X"7480d22e",
        X"84bd3874",
        X"80d22490",
        X"3874bf2e",
        X"9c387480",
        X"d02e81db",
        X"38889239",
        X"7480d32e",
        X"80d93874",
        X"80d72e81",
        X"ca388881",
        X"390282b7",
        X"05330284",
        X"0582b605",
        X"33718280",
        X"29055656",
        X"c9f63f80",
        X"c151c9b0",
        X"3ff4f23f",
        X"fc9e3f83",
        X"c0800883",
        X"c7fc3481",
        X"5283c7fc",
        X"51caca3f",
        X"8151fab1",
        X"3f748e38",
        X"fc823f83",
        X"c0800883",
        X"ca980c87",
        X"39a80b83",
        X"ca980cc9",
        X"bb3f80c1",
        X"51c8f53f",
        X"f4b73f90",
        X"0b83ca93",
        X"33810656",
        X"5674802e",
        X"83389856",
        X"83ca8833",
        X"83ca8933",
        X"71882b07",
        X"56597481",
        X"802e0981",
        X"069c3883",
        X"ca863383",
        X"ca873371",
        X"882b0756",
        X"57ad8075",
        X"278c3875",
        X"81800756",
        X"853975a0",
        X"07567583",
        X"c7fc34ff",
        X"0b83c7fd",
        X"34e00b83",
        X"c7fe3480",
        X"0b83c7ff",
        X"34845283",
        X"c7fc51c9",
        X"bc3f8451",
        X"86b53902",
        X"82b70533",
        X"02840582",
        X"b6053371",
        X"82802905",
        X"565ac8b0",
        X"3f7851ff",
        X"9fb13f83",
        X"c0800880",
        X"2e8a3880",
        X"ce51c7dc",
        X"3f868b39",
        X"80c151c7",
        X"d33fc8c4",
        X"3fc6fd3f",
        X"83caac08",
        X"58837525",
        X"9b3883ca",
        X"883383ca",
        X"89337188",
        X"2b07fc17",
        X"71297a05",
        X"8380055a",
        X"51578d39",
        X"74818029",
        X"18ff8005",
        X"58818057",
        X"80567676",
        X"2e9238c7",
        X"af3f83c0",
        X"800883c7",
        X"fc173481",
        X"1656eb39",
        X"c79e3f83",
        X"c0800881",
        X"ff067753",
        X"83c7fc52",
        X"56f2e23f",
        X"83c08008",
        X"81ff0655",
        X"75752e09",
        X"8106819c",
        X"389451e1",
        X"c53fc798",
        X"3f80c151",
        X"c6d23fc7",
        X"c33f7752",
        X"7851ff9d",
        X"c43f805d",
        X"80d03dfd",
        X"f4055476",
        X"5383c7fc",
        X"527851ff",
        X"9bca3f02",
        X"82b50533",
        X"55815a74",
        X"80d72e09",
        X"810680cc",
        X"38775278",
        X"51ff9d95",
        X"3f80d03d",
        X"fdf00554",
        X"76538e3d",
        X"70537952",
        X"55ff9ccd",
        X"3f805676",
        X"762ea938",
        X"74587770",
        X"81055933",
        X"83c7fc17",
        X"33713270",
        X"30708025",
        X"70307e06",
        X"811b5b5e",
        X"51515155",
        X"75772e09",
        X"8106db38",
        X"82ac51e0",
        X"b93f7980",
        X"2e863880",
        X"c3518439",
        X"80ce51c5",
        X"bf3fc6b0",
        X"3fc4e93f",
        X"83eb3902",
        X"82b70533",
        X"02840582",
        X"b6053371",
        X"82802905",
        X"585a8070",
        X"5c5680e4",
        X"51e0833f",
        X"c5d63f76",
        X"762e0981",
        X"068a3880",
        X"ce51c588",
        X"3f83ba39",
        X"80c151c4",
        X"ff3f83ca",
        X"9408802e",
        X"82d83883",
        X"cab40880",
        X"fc055580",
        X"fd527451",
        X"84a53f83",
        X"c080085a",
        X"768224b2",
        X"38ff1770",
        X"872b83ff",
        X"ff800680",
        X"fdcc0583",
        X"c7fc5957",
        X"55818055",
        X"75708105",
        X"57337770",
        X"81055934",
        X"ff157081",
        X"ff065155",
        X"74ea3882",
        X"87397682",
        X"e82e81a5",
        X"387682e9",
        X"2e098106",
        X"81ac3875",
        X"765a5877",
        X"87327030",
        X"70720780",
        X"257a8a32",
        X"70307072",
        X"07802573",
        X"0753545a",
        X"51575575",
        X"802e9738",
        X"78782692",
        X"38a00b83",
        X"c7fc1a34",
        X"81197081",
        X"ff065a55",
        X"eb398118",
        X"7081ff06",
        X"59558a78",
        X"27ffbc38",
        X"8f5883c7",
        X"f7183383",
        X"c7fc1934",
        X"ff187081",
        X"ff065955",
        X"778426ea",
        X"38905880",
        X"0b83c7fc",
        X"19348118",
        X"7081ff06",
        X"70982b52",
        X"59557480",
        X"25e93880",
        X"c6557985",
        X"8f248438",
        X"80c25574",
        X"83c7fc34",
        X"80f10b83",
        X"c7ff3481",
        X"0b83c880",
        X"347983c7",
        X"fd347988",
        X"2c557483",
        X"c7fe3480",
        X"cb3982f0",
        X"772580c4",
        X"387680fd",
        X"29fd97d3",
        X"05527851",
        X"ff99d63f",
        X"80d03dfd",
        X"ec055480",
        X"fd5383c7",
        X"fc527851",
        X"ff998e3f",
        X"7a811858",
        X"587780fc",
        X"24833875",
        X"5776882c",
        X"557483c8",
        X"f9347683",
        X"c8fa3477",
        X"83c8fb34",
        X"81805680",
        X"cc3983ca",
        X"ac085883",
        X"77259b38",
        X"83ca8833",
        X"83ca8933",
        X"71882b07",
        X"fc197129",
        X"7a058380",
        X"055a575a",
        X"8d397681",
        X"802918ff",
        X"80055881",
        X"80567752",
        X"7851ff98",
        X"e43f80d0",
        X"3dfdec05",
        X"54755383",
        X"c7fc5278",
        X"51ff989d",
        X"3f7551f2",
        X"ec3fc2c0",
        X"3fc0f93f",
        X"8b3983c9",
        X"fc088105",
        X"83c9fc0c",
        X"80d03d0d",
        X"04f6c03f",
        X"fc39dc89",
        X"3f04803d",
        X"0ddc823f",
        X"83c08008",
        X"842980ff",
        X"a0057008",
        X"83c0800c",
        X"51823d0d",
        X"04fc3d0d",
        X"76785354",
        X"81538055",
        X"87397110",
        X"73105452",
        X"73722651",
        X"72802ea7",
        X"3870802e",
        X"86387180",
        X"25e83872",
        X"802e9838",
        X"71742689",
        X"38737231",
        X"75740756",
        X"5472812a",
        X"72812a53",
        X"53e53973",
        X"51788338",
        X"74517083",
        X"c0800c86",
        X"3d0d04fe",
        X"3d0d8053",
        X"75527451",
        X"ffa33f84",
        X"3d0d04fe",
        X"3d0d8153",
        X"75527451",
        X"ff933f84",
        X"3d0d04fb",
        X"3d0d7779",
        X"55558056",
        X"74762586",
        X"38743055",
        X"81567380",
        X"25883873",
        X"30768132",
        X"57548053",
        X"73527451",
        X"fee73f83",
        X"c0800854",
        X"75802e87",
        X"3883c080",
        X"08305473",
        X"83c0800c",
        X"873d0d04",
        X"fa3d0d78",
        X"7a575580",
        X"57747725",
        X"86387430",
        X"55815775",
        X"9f2c5481",
        X"53757432",
        X"74315274",
        X"51feaa3f",
        X"83c08008",
        X"5476802e",
        X"873883c0",
        X"80083054",
        X"7383c080",
        X"0c883d0d",
        X"04fd3d0d",
        X"75548074",
        X"0c800b84",
        X"150c800b",
        X"88150c80",
        X"0b8c150c",
        X"87a68033",
        X"7081ff06",
        X"7071842a",
        X"06515151",
        X"d9be3f70",
        X"812a8132",
        X"71813271",
        X"81067181",
        X"06318417",
        X"0c535370",
        X"832a8132",
        X"71822a81",
        X"32708106",
        X"72713177",
        X"0c515252",
        X"87a09033",
        X"87a09133",
        X"7081ff06",
        X"70730681",
        X"32810688",
        X"180c5152",
        X"5283c080",
        X"08802e80",
        X"c23883c0",
        X"8008812a",
        X"70810683",
        X"c0800881",
        X"06318416",
        X"0c5183c0",
        X"8008832a",
        X"83c08008",
        X"822a7181",
        X"06718106",
        X"31760c52",
        X"5283c080",
        X"08842a81",
        X"0688150c",
        X"83c08008",
        X"852a8106",
        X"8c150c85",
        X"3d0d04fe",
        X"3d0d7476",
        X"54527151",
        X"febb3fd7",
        X"f53f83c0",
        X"8008802e",
        X"8938810b",
        X"8c130c80",
        X"d0397281",
        X"2ea73881",
        X"73268d38",
        X"72822ead",
        X"3872832e",
        X"a138d339",
        X"7108cf38",
        X"841208ca",
        X"38881208",
        X"c5388c12",
        X"08c038a5",
        X"39881208",
        X"812e9e38",
        X"91398812",
        X"08812e95",
        X"38710891",
        X"38841208",
        X"8c388c12",
        X"08812e09",
        X"8106ff9a",
        X"38843d0d",
        X"04000000",
        X"00ffffff",
        X"ff00ffff",
        X"ffff00ff",
        X"ffffff00",
        X"809a9041",
        X"8e418f80",
        X"45454549",
        X"49498e8f",
        X"9092924f",
        X"994f5555",
        X"59999a9b",
        X"9c9d9e9f",
        X"41494f55",
        X"a5a5a6a7",
        X"a8a9aaab",
        X"ac21aeaf",
        X"b0b1b2b3",
        X"b4b5b6b7",
        X"b8b9babb",
        X"bcbdbebf",
        X"c0c1c2c3",
        X"c4c5c6c7",
        X"c8c9cacb",
        X"cccdcecf",
        X"d0d1d2d3",
        X"d4d5d6d7",
        X"d8d9dadb",
        X"dcdddedf",
        X"e0e1e2e3",
        X"e4e5e6e7",
        X"e8e9eaeb",
        X"ecedeeef",
        X"f0f1f2f3",
        X"f4f5f6f7",
        X"f8f9fafb",
        X"fcfdfeff",
        X"00000000",
        X"00002bcb",
        X"00002bf1",
        X"00002bf1",
        X"00002bf1",
        X"00002bf1",
        X"00002c62",
        X"00002cb3",
        X"2e2e0000",
        X"41545200",
        X"58464400",
        X"58455800",
        X"43686f6f",
        X"73652000",
        X"66696c65",
        X"00000000",
        X"4449523a",
        X"00000000",
        X"44495200",
        X"25732025",
        X"73000000",
        X"20000000",
        X"25303278",
        X"00000000",
        X"53650000",
        X"7474696e",
        X"67730000",
        X"526f6d3a",
        X"25730000",
        X"44726976",
        X"65202564",
        X"3a257320",
        X"25730000",
        X"4e4f4e45",
        X"00000000",
        X"43617274",
        X"3a202573",
        X"00000000",
        X"45786974",
        X"00000000",
        X"61746172",
        X"69626173",
        X"2e726f6d",
        X"00000000",
        X"61746172",
        X"69786c2e",
        X"726f6d00",
        X"61746172",
        X"696f7362",
        X"2e726f6d",
        X"00000000",
        X"66726565",
        X"7a65722e",
        X"726f6d00",
        X"524f4d00",
        X"42494e00",
        X"43415200",
        X"4d454d00",
        X"5374616e",
        X"64617264",
        X"00000000",
        X"46617374",
        X"28362900",
        X"46617374",
        X"28352900",
        X"46617374",
        X"28342900",
        X"46617374",
        X"28332900",
        X"46617374",
        X"28322900",
        X"46617374",
        X"28312900",
        X"46617374",
        X"28302900",
        X"00000000",
        X"00000000",
        X"01010008",
        X"02210010",
        X"080d0040",
        X"090a0040",
        X"0a090040",
        X"0b080040",
        X"0c300020",
        X"0d310040",
        X"0e320080",
        X"0f040010",
        X"110c0080",
        X"17330100",
        X"18340200",
        X"1a280010",
        X"1b290020",
        X"1c2a0040",
        X"1d2b0080",
        X"1e2c0100",
        X"1f2d0200",
        X"21380020",
        X"22390040",
        X"233a0080",
        X"243b0100",
        X"253c0200",
        X"28230010",
        X"29020080",
        X"2a030400",
        X"38240200",
        X"00000000",
        X"70704740",
        X"2c704268",
        X"2c020202",
        X"02020202",
        X"02020202",
        X"02020202",
        X"02020202",
        X"02020241",
        X"00060000",
        X"72025f07",
        X"f807a900",
        X"8d04038d",
        X"4402a907",
        X"8d0503a9",
        X"708d0a03",
        X"a9018d0b",
        X"03850960",
        X"7d8a4820",
        X"53e488d0",
        X"fa68aa8c",
        X"8e07ad7d",
        X"07ee8e07",
        X"60a9938d",
        X"e202a907",
        X"8de302a2",
        X"0220da07",
        X"954320da",
        X"07954435",
        X"43c9fff0",
        X"f0caca10",
        X"ec3006e6",
        X"45d002e6",
        X"4620da07",
        X"a2018144",
        X"b545d543",
        X"d0edca10",
        X"f720d207",
        X"4c9407a9",
        X"038d0fd2",
        X"6ce202ad",
        X"8e07cd7f",
        X"07d0abee",
        X"0a03d003",
        X"ee0b03ad",
        X"7d070d7e",
        X"07d08e20",
        X"d2076ce0",
        X"0220da07",
        X"8de00220",
        X"da078de1",
        X"022de002",
        X"c9fff0ed",
        X"a9008d8e",
        X"07f08200",
        X"00000028",
        X"00000006",
        X"00000005",
        X"00000004",
        X"00000003",
        X"00000002",
        X"00000001",
        X"00000000",
        X"00003de8",
        X"00003df4",
        X"00003dfc",
        X"00003e04",
        X"00003e0c",
        X"00003e14",
        X"00003e1c",
        X"00003e24",
        X"2f617461",
        X"72693830",
        X"302f726f",
        X"6d000000",
        X"2f617461",
        X"72693830",
        X"302f7573",
        X"65720000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000"

);

signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
