
--
--ROMsUsingBlockRAMResources.
--VHDLcodeforaROMwithregisteredoutput(template2)
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity zpu_rom is
port(
        clock:in std_logic;
        address:in std_logic_vector(11 downto 0);
        q:out std_logic_vector(31 downto 0)
);
end zpu_rom;

architecture syn of zpu_rom is
        type rom_type is array(0 to 4095) of std_logic_vector(31 downto 0);
        signal ROM:rom_type:=
(
        X"0b0b0b89",
        X"ad040b0b",
        X"0b0b0b0b",
        X"0b0b0b0b",
        X"0b0b0b0b",
        X"0b0b0b0b",
        X"0b0b0b0b",
        X"0b0b0b0b",
        X"0b0b0b0b",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"71fd0608",
        X"72830609",
        X"81058205",
        X"832b2a83",
        X"ffff0652",
        X"04000000",
        X"00000000",
        X"00000000",
        X"71fd0608",
        X"83ffff73",
        X"83060981",
        X"05820583",
        X"2b2b0906",
        X"7383ffff",
        X"0b0b0b0b",
        X"83a70400",
        X"72098105",
        X"72057373",
        X"09060906",
        X"73097306",
        X"070a8106",
        X"53510400",
        X"00000000",
        X"00000000",
        X"72722473",
        X"732e0753",
        X"51040000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"71737109",
        X"71068106",
        X"30720a10",
        X"0a720a10",
        X"0a31050a",
        X"81065151",
        X"53510400",
        X"00000000",
        X"72722673",
        X"732e0753",
        X"51040000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"0b0b0b88",
        X"bc040000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"720a722b",
        X"0a535104",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"72729f06",
        X"0981050b",
        X"0b0b889f",
        X"05040000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"72722aff",
        X"739f062a",
        X"0974090a",
        X"8106ff05",
        X"06075351",
        X"04000000",
        X"00000000",
        X"00000000",
        X"71715351",
        X"020d0406",
        X"73830609",
        X"81058205",
        X"832b0b2b",
        X"0772fc06",
        X"0c515104",
        X"00000000",
        X"72098105",
        X"72050970",
        X"81050906",
        X"0a810653",
        X"51040000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"72098105",
        X"72050970",
        X"81050906",
        X"0a098106",
        X"53510400",
        X"00000000",
        X"00000000",
        X"00000000",
        X"71098105",
        X"52040000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"72720981",
        X"05055351",
        X"04000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"72097206",
        X"73730906",
        X"07535104",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"71fc0608",
        X"72830609",
        X"81058305",
        X"1010102a",
        X"81ff0652",
        X"04000000",
        X"00000000",
        X"00000000",
        X"71fc0608",
        X"0b0b80e9",
        X"80738306",
        X"10100508",
        X"060b0b0b",
        X"88a20400",
        X"00000000",
        X"00000000",
        X"0b0b0b88",
        X"ff040000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"0b0b0b88",
        X"d8040000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"72097081",
        X"0509060a",
        X"8106ff05",
        X"70547106",
        X"73097274",
        X"05ff0506",
        X"07515151",
        X"04000000",
        X"72097081",
        X"0509060a",
        X"098106ff",
        X"05705471",
        X"06730972",
        X"7405ff05",
        X"06075151",
        X"51040000",
        X"05ff0504",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"810b80ec",
        X"d80c5104",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00007181",
        X"05520400",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000284",
        X"05721010",
        X"05520400",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00007171",
        X"05ff0571",
        X"5351020d",
        X"04000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"10101010",
        X"10101010",
        X"10101010",
        X"10101010",
        X"10101010",
        X"10101010",
        X"10101010",
        X"10101053",
        X"51047381",
        X"ff067383",
        X"06098105",
        X"83051010",
        X"102b0772",
        X"fc060c51",
        X"51043c04",
        X"72728072",
        X"8106ff05",
        X"09720605",
        X"71105272",
        X"0a100a53",
        X"72ed3851",
        X"51535104",
        X"83e08008",
        X"83e08408",
        X"83e08808",
        X"757580e7",
        X"9b2d5050",
        X"83e08008",
        X"5683e088",
        X"0c83e084",
        X"0c83e080",
        X"0c510483",
        X"e0800883",
        X"e0840883",
        X"e0880875",
        X"7580e6da",
        X"2d505083",
        X"e0800856",
        X"83e0880c",
        X"83e0840c",
        X"83e0800c",
        X"51040000",
        X"800489aa",
        X"0489aa0b",
        X"80e0a704",
        X"fd3d0d75",
        X"705254af",
        X"bb3f83e0",
        X"80081453",
        X"72742e92",
        X"38ff1370",
        X"33535371",
        X"af2e0981",
        X"06ee3881",
        X"13537283",
        X"e0800c85",
        X"3d0d04fd",
        X"3d0d7577",
        X"70535454",
        X"c73f83e0",
        X"8008732e",
        X"a13883e0",
        X"80087331",
        X"52ff1252",
        X"71ff2e8f",
        X"38727081",
        X"05543374",
        X"70810556",
        X"34eb39ff",
        X"14548074",
        X"34853d0d",
        X"04803d0d",
        X"7251ff90",
        X"3f823d0d",
        X"047183e0",
        X"800c0480",
        X"3d0d7251",
        X"80713481",
        X"0bbc120c",
        X"800b80c0",
        X"120c823d",
        X"0d04800b",
        X"83e2c008",
        X"248a38b6",
        X"8c3fff0b",
        X"83e2c00c",
        X"800b83e0",
        X"800c04ff",
        X"3d0d7352",
        X"83e09c08",
        X"722e8d38",
        X"d93f7151",
        X"96a03f71",
        X"83e09c0c",
        X"833d0d04",
        X"f43d0d7e",
        X"60625c5a",
        X"55805681",
        X"54bc1508",
        X"762e0981",
        X"06819138",
        X"7451c83f",
        X"7958757a",
        X"2580f738",
        X"83e2f008",
        X"70892a57",
        X"83ff0678",
        X"84807231",
        X"56565773",
        X"78258338",
        X"73557583",
        X"e2c0082e",
        X"8438ff82",
        X"3f83e2c0",
        X"088025a6",
        X"3875892b",
        X"5198dc3f",
        X"83e2f008",
        X"8f3dfc11",
        X"555c5481",
        X"52f81b51",
        X"96c63f76",
        X"1483e2f0",
        X"0c7583e2",
        X"c00c7453",
        X"76527851",
        X"b4b63f83",
        X"e0800883",
        X"e2f00816",
        X"83e2f00c",
        X"78763176",
        X"1b5b5956",
        X"778024ff",
        X"8b38617a",
        X"710c5475",
        X"5475802e",
        X"83388154",
        X"7383e080",
        X"0c8e3d0d",
        X"04fc3d0d",
        X"fe943f76",
        X"51fea83f",
        X"863dfc05",
        X"53785277",
        X"5195e93f",
        X"7975710c",
        X"5483e080",
        X"085483e0",
        X"8008802e",
        X"83388154",
        X"7383e080",
        X"0c863d0d",
        X"04fe3d0d",
        X"7583e2c0",
        X"08535380",
        X"72248938",
        X"71732e84",
        X"38fdcf3f",
        X"7451fde3",
        X"3f725197",
        X"ae3f83e0",
        X"80085283",
        X"e0800880",
        X"2e833881",
        X"527183e0",
        X"800c843d",
        X"0d04803d",
        X"0d7280c0",
        X"110883e0",
        X"800c5182",
        X"3d0d0480",
        X"3d0d72bc",
        X"110883e0",
        X"800c5182",
        X"3d0d0480",
        X"c40b83e0",
        X"800c04fd",
        X"3d0d7577",
        X"71547053",
        X"5553ab8c",
        X"3f82c813",
        X"08bc150c",
        X"82c01308",
        X"80c0150c",
        X"fce43f73",
        X"5193ab3f",
        X"7383e09c",
        X"0c83e080",
        X"085383e0",
        X"8008802e",
        X"83388153",
        X"7283e080",
        X"0c853d0d",
        X"04fd3d0d",
        X"75775553",
        X"fcb83f72",
        X"802ea538",
        X"bc130852",
        X"7351aa96",
        X"3f83e080",
        X"088f3877",
        X"527251ff",
        X"9a3f83e0",
        X"8008538a",
        X"3982cc13",
        X"0853d839",
        X"81537283",
        X"e0800c85",
        X"3d0d04fe",
        X"3d0dff0b",
        X"83e2c00c",
        X"7483e0a0",
        X"0c7583e2",
        X"bc0cb0ea",
        X"3f83e080",
        X"0881ff06",
        X"52815371",
        X"993883e2",
        X"d8518e94",
        X"3f83e080",
        X"085283e0",
        X"8008802e",
        X"83387252",
        X"71537283",
        X"e0800c84",
        X"3d0d04fa",
        X"3d0d787a",
        X"82c41208",
        X"82c41208",
        X"70722459",
        X"56565757",
        X"73732e09",
        X"81069138",
        X"80c01652",
        X"80c01751",
        X"a8873f83",
        X"e0800855",
        X"7483e080",
        X"0c883d0d",
        X"04f63d0d",
        X"7c5b807b",
        X"715c5457",
        X"7a772e8c",
        X"38811a82",
        X"cc140854",
        X"5a72f638",
        X"805980d9",
        X"397a5481",
        X"5780707b",
        X"7b315a57",
        X"55ff1853",
        X"74732580",
        X"c13882cc",
        X"14085273",
        X"51ff8c3f",
        X"800b83e0",
        X"800825a1",
        X"3882cc14",
        X"0882cc11",
        X"0882cc16",
        X"0c7482cc",
        X"120c5375",
        X"802e8638",
        X"7282cc17",
        X"0c725480",
        X"577382cc",
        X"15088117",
        X"575556ff",
        X"b8398119",
        X"59800bff",
        X"1b545478",
        X"73258338",
        X"81547681",
        X"32707506",
        X"515372ff",
        X"90388c3d",
        X"0d04f73d",
        X"0d7b7d5a",
        X"5a82d052",
        X"83e2bc08",
        X"5180d5d6",
        X"3f83e080",
        X"0857f9da",
        X"3f795283",
        X"e2c45195",
        X"b73f83e0",
        X"80085480",
        X"5383e080",
        X"08732e09",
        X"81068283",
        X"3883e0a0",
        X"080b0b80",
        X"eacc5370",
        X"5256a7c4",
        X"3f0b0b80",
        X"eacc5280",
        X"c01651a7",
        X"b73f75bc",
        X"170c7382",
        X"c0170c81",
        X"0b82c417",
        X"0c810b82",
        X"c8170c73",
        X"82cc170c",
        X"ff1782d0",
        X"17555781",
        X"913983e0",
        X"ac337082",
        X"2a708106",
        X"51545572",
        X"81803874",
        X"812a8106",
        X"587780f6",
        X"3874842a",
        X"810682c4",
        X"150c83e0",
        X"ac338106",
        X"82c8150c",
        X"79527351",
        X"a6de3f73",
        X"51a6f53f",
        X"83e08008",
        X"1453af73",
        X"70810555",
        X"3472bc15",
        X"0c83e0ad",
        X"527251a6",
        X"bf3f83e0",
        X"a40882c0",
        X"150c83e0",
        X"ba5280c0",
        X"1451a6ac",
        X"3f78802e",
        X"8d387351",
        X"782d83e0",
        X"8008802e",
        X"99387782",
        X"cc150c75",
        X"802e8638",
        X"7382cc17",
        X"0c7382d0",
        X"15ff1959",
        X"55567680",
        X"2e9b3883",
        X"e0a45283",
        X"e2c45194",
        X"ad3f83e0",
        X"80088a38",
        X"83e0ad33",
        X"5372fed2",
        X"3878802e",
        X"893883e0",
        X"a00851fc",
        X"b83f83e0",
        X"a0085372",
        X"83e0800c",
        X"8b3d0d04",
        X"ff3d0d80",
        X"527351fd",
        X"b53f833d",
        X"0d04f03d",
        X"0d627052",
        X"54f6893f",
        X"83e08008",
        X"7453873d",
        X"70535555",
        X"f6a93ff7",
        X"893f7351",
        X"d33f6353",
        X"745283e0",
        X"800851fa",
        X"b83f923d",
        X"0d047183",
        X"e0800c04",
        X"80c01283",
        X"e0800c04",
        X"803d0d72",
        X"82c01108",
        X"83e0800c",
        X"51823d0d",
        X"04803d0d",
        X"7282cc11",
        X"0883e080",
        X"0c51823d",
        X"0d04803d",
        X"0d7282c4",
        X"110883e0",
        X"800c5182",
        X"3d0d04f9",
        X"3d0d7983",
        X"e0900857",
        X"57817727",
        X"81963876",
        X"88170827",
        X"818e3875",
        X"33557482",
        X"2e893874",
        X"832eb338",
        X"80fe3974",
        X"54761083",
        X"fe065376",
        X"882a8c17",
        X"08055289",
        X"3dfc0551",
        X"ab983f83",
        X"e0800880",
        X"df38029d",
        X"0533893d",
        X"3371882b",
        X"07565680",
        X"d1398454",
        X"76822b83",
        X"fc065376",
        X"872a8c17",
        X"08055289",
        X"3dfc0551",
        X"aae83f83",
        X"e08008b0",
        X"38029f05",
        X"33028405",
        X"9e053371",
        X"982b7190",
        X"2b07028c",
        X"059d0533",
        X"70882b72",
        X"078d3d33",
        X"7180ffff",
        X"fe800607",
        X"51525357",
        X"58568339",
        X"81557483",
        X"e0800c89",
        X"3d0d04fb",
        X"3d0d83e0",
        X"9008fe19",
        X"881208fe",
        X"05555654",
        X"80567473",
        X"278d3882",
        X"14337571",
        X"29941608",
        X"05575375",
        X"83e0800c",
        X"873d0d04",
        X"fc3d0d76",
        X"52800b83",
        X"e0900870",
        X"33515253",
        X"70832e09",
        X"81069138",
        X"95123394",
        X"13337198",
        X"2b71902b",
        X"07555551",
        X"9b12339a",
        X"13337188",
        X"2b077407",
        X"83e0800c",
        X"55863d0d",
        X"04fc3d0d",
        X"7683e090",
        X"08555580",
        X"75238815",
        X"08537281",
        X"2e883888",
        X"14087326",
        X"85388152",
        X"b2397290",
        X"38733352",
        X"71832e09",
        X"81068538",
        X"90140853",
        X"728c160c",
        X"72802e8d",
        X"387251fe",
        X"d63f83e0",
        X"80085285",
        X"39901408",
        X"52719016",
        X"0c805271",
        X"83e0800c",
        X"863d0d04",
        X"fa3d0d78",
        X"83e09008",
        X"71228105",
        X"7083ffff",
        X"06575457",
        X"5573802e",
        X"88389015",
        X"08537286",
        X"38835280",
        X"e739738f",
        X"06527180",
        X"da388113",
        X"90160c8c",
        X"15085372",
        X"9038830b",
        X"84172257",
        X"52737627",
        X"80c638bf",
        X"39821633",
        X"ff057484",
        X"2a065271",
        X"b2387251",
        X"fcb13f81",
        X"527183e0",
        X"800827a8",
        X"38835283",
        X"e0800888",
        X"1708279c",
        X"3883e080",
        X"088c160c",
        X"83e08008",
        X"51fdbc3f",
        X"83e08008",
        X"90160c73",
        X"75238052",
        X"7183e080",
        X"0c883d0d",
        X"04f23d0d",
        X"60626458",
        X"5e5b7533",
        X"5574a02e",
        X"09810688",
        X"38811670",
        X"4456ef39",
        X"62703356",
        X"5674af2e",
        X"09810684",
        X"38811643",
        X"800b881c",
        X"0c627033",
        X"5155749f",
        X"2691387a",
        X"51fdd23f",
        X"83e08008",
        X"56807d34",
        X"83813993",
        X"3d841c08",
        X"7058595f",
        X"8a55a076",
        X"70810558",
        X"34ff1555",
        X"74ff2e09",
        X"8106ef38",
        X"80705a5c",
        X"887f085f",
        X"5a7b811d",
        X"7081ff06",
        X"60137033",
        X"70af3270",
        X"30a07327",
        X"71802507",
        X"5151525b",
        X"535e5755",
        X"7480e738",
        X"76ae2e09",
        X"81068338",
        X"8155787a",
        X"27750755",
        X"74802e9f",
        X"38798832",
        X"703078ae",
        X"32703070",
        X"73079f2a",
        X"53515751",
        X"5675bb38",
        X"88598b5a",
        X"ffab3976",
        X"982b5574",
        X"80258738",
        X"80e89017",
        X"3357ff9f",
        X"17557499",
        X"268938e0",
        X"177081ff",
        X"06585578",
        X"811a7081",
        X"ff067a13",
        X"535b5755",
        X"767534fe",
        X"f8397b1e",
        X"7f0c8055",
        X"76a02683",
        X"38815574",
        X"8b19347a",
        X"51fc823f",
        X"83e08008",
        X"80f538a0",
        X"547a2270",
        X"852b83e0",
        X"06545590",
        X"1b08527c",
        X"51a5a33f",
        X"83e08008",
        X"5783e080",
        X"08818138",
        X"7c335574",
        X"802e80f4",
        X"388b1d33",
        X"70832a70",
        X"81065156",
        X"5674b438",
        X"8b7d841d",
        X"0883e080",
        X"08595b5b",
        X"58ff1858",
        X"77ff2e9a",
        X"38797081",
        X"055b3379",
        X"7081055b",
        X"33717131",
        X"52565675",
        X"802ee238",
        X"86397580",
        X"2e96387a",
        X"51fbe53f",
        X"ff863983",
        X"e0800856",
        X"83e08008",
        X"b6388339",
        X"7656841b",
        X"088b1133",
        X"515574a7",
        X"388b1d33",
        X"70842a70",
        X"81065156",
        X"56748938",
        X"83569439",
        X"81569039",
        X"7c51fa94",
        X"3f83e080",
        X"08881c0c",
        X"fd813975",
        X"83e0800c",
        X"903d0d04",
        X"f83d0d7a",
        X"7c595782",
        X"5483fe53",
        X"77527651",
        X"a3e83f83",
        X"5683e080",
        X"0880ec38",
        X"81173377",
        X"3371882b",
        X"07565682",
        X"567482d4",
        X"d52e0981",
        X"0680d438",
        X"7554b653",
        X"77527651",
        X"a3bc3f83",
        X"e0800898",
        X"38811733",
        X"77337188",
        X"2b0783e0",
        X"80085256",
        X"56748182",
        X"c62eac38",
        X"825480d2",
        X"53775276",
        X"51a3933f",
        X"83e08008",
        X"98388117",
        X"33773371",
        X"882b0783",
        X"e0800852",
        X"56567481",
        X"82c62e83",
        X"38815675",
        X"83e0800c",
        X"8a3d0d04",
        X"eb3d0d67",
        X"5a800b83",
        X"e0900ca2",
        X"b53f83e0",
        X"80088106",
        X"55825674",
        X"83ef3874",
        X"75538f3d",
        X"70535759",
        X"feca3f83",
        X"e0800881",
        X"ff065776",
        X"812e0981",
        X"0680d438",
        X"905483be",
        X"53745275",
        X"51a2a73f",
        X"83e08008",
        X"80c9388f",
        X"3d335574",
        X"802e80c9",
        X"3802bf05",
        X"33028405",
        X"be053371",
        X"982b7190",
        X"2b07028c",
        X"05bd0533",
        X"70882b72",
        X"07953d33",
        X"71077058",
        X"7b575e52",
        X"5e575957",
        X"fdee3f83",
        X"e0800881",
        X"ff065776",
        X"832e0981",
        X"06863881",
        X"5682f239",
        X"76802e86",
        X"38865682",
        X"e839a454",
        X"8d537852",
        X"7551a1be",
        X"3f815683",
        X"e0800882",
        X"d43802be",
        X"05330284",
        X"05bd0533",
        X"71882b07",
        X"595d77ab",
        X"380280ce",
        X"05330284",
        X"0580cd05",
        X"3371982b",
        X"71902b07",
        X"973d3370",
        X"882b7207",
        X"02940580",
        X"cb053371",
        X"0754525e",
        X"57595602",
        X"b7053378",
        X"71290288",
        X"05b60533",
        X"028c05b5",
        X"05337188",
        X"2b07701d",
        X"707f8c05",
        X"0c5f5957",
        X"595d8e3d",
        X"33821b34",
        X"02b90533",
        X"903d3371",
        X"882b075a",
        X"5c78841b",
        X"2302bb05",
        X"33028405",
        X"ba053371",
        X"882b0756",
        X"5c74ab38",
        X"0280ca05",
        X"33028405",
        X"80c90533",
        X"71982b71",
        X"902b0796",
        X"3d337088",
        X"2b720702",
        X"940580c7",
        X"05337107",
        X"51525357",
        X"5e5c7476",
        X"31783179",
        X"842a903d",
        X"33547171",
        X"31535656",
        X"80c6bb3f",
        X"83e08008",
        X"82057088",
        X"1c0c83e0",
        X"8008e08a",
        X"05565674",
        X"83dffe26",
        X"83388257",
        X"83fff676",
        X"27853883",
        X"57893986",
        X"5676802e",
        X"80db3876",
        X"7a347683",
        X"2e098106",
        X"b0380280",
        X"d6053302",
        X"840580d5",
        X"05337198",
        X"2b71902b",
        X"07993d33",
        X"70882b72",
        X"07029405",
        X"80d30533",
        X"71077f90",
        X"050c525e",
        X"57585686",
        X"39771b90",
        X"1b0c841a",
        X"228c1b08",
        X"1971842a",
        X"05941c0c",
        X"5d800b81",
        X"1b347983",
        X"e0900c80",
        X"567583e0",
        X"800c973d",
        X"0d04e93d",
        X"0d83e090",
        X"08568554",
        X"75802e81",
        X"8238800b",
        X"81173499",
        X"3de01146",
        X"6a548a3d",
        X"705458ec",
        X"0551f6e5",
        X"3f83e080",
        X"085483e0",
        X"800880df",
        X"38893d33",
        X"5473802e",
        X"913802ab",
        X"05337084",
        X"2a810651",
        X"5574802e",
        X"86388354",
        X"80c13976",
        X"51f4893f",
        X"83e08008",
        X"a0170c02",
        X"bf053302",
        X"8405be05",
        X"3371982b",
        X"71902b07",
        X"028c05bd",
        X"05337088",
        X"2b720795",
        X"3d337107",
        X"9c1c0c52",
        X"78981b0c",
        X"53565957",
        X"810b8117",
        X"34745473",
        X"83e0800c",
        X"993d0d04",
        X"f53d0d7d",
        X"7f617283",
        X"e090085a",
        X"5d5d595c",
        X"807b0c85",
        X"5775802e",
        X"81e03881",
        X"16338106",
        X"55845774",
        X"802e81d2",
        X"38913974",
        X"81173486",
        X"39800b81",
        X"17348157",
        X"81c0399c",
        X"16089817",
        X"08315574",
        X"78278338",
        X"74587780",
        X"2e81a938",
        X"98160870",
        X"83ff0656",
        X"577480cf",
        X"38821633",
        X"ff057789",
        X"2a067081",
        X"ff065a55",
        X"78a03876",
        X"8738a016",
        X"08558d39",
        X"a4160851",
        X"f0e93f83",
        X"e0800855",
        X"817527ff",
        X"a83874a4",
        X"170ca416",
        X"0851f283",
        X"3f83e080",
        X"085583e0",
        X"8008802e",
        X"ff893883",
        X"e0800819",
        X"a8170c98",
        X"160883ff",
        X"06848071",
        X"31515577",
        X"75278338",
        X"77557483",
        X"ffff0654",
        X"98160883",
        X"ff0653a8",
        X"16085279",
        X"577b8338",
        X"7b577651",
        X"9be43f83",
        X"e08008fe",
        X"d0389816",
        X"08159817",
        X"0c741a78",
        X"76317c08",
        X"177d0c59",
        X"5afed339",
        X"80577683",
        X"e0800c8d",
        X"3d0d04fa",
        X"3d0d7883",
        X"e0900855",
        X"56855573",
        X"802e81e3",
        X"38811433",
        X"81065384",
        X"5572802e",
        X"81d5389c",
        X"14085372",
        X"76278338",
        X"72569814",
        X"0857800b",
        X"98150c75",
        X"802e81b9",
        X"38821433",
        X"70892b56",
        X"5376802e",
        X"b7387452",
        X"ff165180",
        X"c1bc3f83",
        X"e08008ff",
        X"18765470",
        X"53585380",
        X"c1ac3f83",
        X"e0800873",
        X"26963874",
        X"30707806",
        X"7098170c",
        X"777131a4",
        X"17085258",
        X"51538939",
        X"a0140870",
        X"a4160c53",
        X"747627b9",
        X"387251ee",
        X"d63f83e0",
        X"80085381",
        X"0b83e080",
        X"08278b38",
        X"88140883",
        X"e0800826",
        X"8838800b",
        X"811534b0",
        X"3983e080",
        X"08a4150c",
        X"98140815",
        X"98150c75",
        X"753156c4",
        X"39981408",
        X"16709816",
        X"0c735256",
        X"efc53f83",
        X"e080088c",
        X"3883e080",
        X"08811534",
        X"81559439",
        X"821433ff",
        X"0576892a",
        X"0683e080",
        X"0805a815",
        X"0c805574",
        X"83e0800c",
        X"883d0d04",
        X"ef3d0d63",
        X"56855583",
        X"e0900880",
        X"2e80d238",
        X"933df405",
        X"84170c64",
        X"53883d70",
        X"53765257",
        X"f1cf3f83",
        X"e0800855",
        X"83e08008",
        X"b438883d",
        X"33547380",
        X"2ea13802",
        X"a7053370",
        X"842a7081",
        X"06515555",
        X"83557380",
        X"2e973876",
        X"51eef53f",
        X"83e08008",
        X"88170c75",
        X"51efa63f",
        X"83e08008",
        X"557483e0",
        X"800c933d",
        X"0d04e43d",
        X"0d6ea13d",
        X"08405e85",
        X"5683e090",
        X"08802e84",
        X"85389e3d",
        X"f405841f",
        X"0c7e9838",
        X"7d51eef5",
        X"3f83e080",
        X"085683ee",
        X"39814181",
        X"f6398341",
        X"81f13993",
        X"3d7f9605",
        X"4159807f",
        X"8295055e",
        X"56756081",
        X"ff053483",
        X"41901e08",
        X"762e81d3",
        X"38a0547d",
        X"2270852b",
        X"83e00654",
        X"58901e08",
        X"52785197",
        X"ed3f83e0",
        X"80084183",
        X"e08008ff",
        X"b8387833",
        X"5c7b802e",
        X"ffb4388b",
        X"193370bf",
        X"06718106",
        X"52435574",
        X"802e80de",
        X"387b81bf",
        X"0655748f",
        X"2480d338",
        X"9a193355",
        X"7480cb38",
        X"f31d7058",
        X"5d815675",
        X"8b2e0981",
        X"0685388e",
        X"568b3975",
        X"9a2e0981",
        X"0683389c",
        X"56781670",
        X"70810552",
        X"33713381",
        X"1a821a5f",
        X"5b525b55",
        X"74863879",
        X"77348539",
        X"80df7734",
        X"777b5757",
        X"7aa02e09",
        X"8106c038",
        X"81567b81",
        X"e5327030",
        X"709f2a51",
        X"51557bae",
        X"2e933874",
        X"802e8e38",
        X"61832a70",
        X"81065155",
        X"74802e97",
        X"387d51ed",
        X"df3f83e0",
        X"80084183",
        X"e0800887",
        X"38901e08",
        X"feaf3880",
        X"60347580",
        X"2e88387c",
        X"527f518f",
        X"933f6080",
        X"2e863880",
        X"0b901f0c",
        X"60566083",
        X"2e853860",
        X"81d03889",
        X"1f57901e",
        X"08802e81",
        X"a8388056",
        X"78167033",
        X"515574a0",
        X"2ea03874",
        X"852e0981",
        X"06843881",
        X"e5557477",
        X"70810559",
        X"34811670",
        X"81ff0657",
        X"55877627",
        X"d7388819",
        X"335574a0",
        X"2ea938ae",
        X"77708105",
        X"59348856",
        X"78167033",
        X"515574a0",
        X"2e953874",
        X"77708105",
        X"59348116",
        X"7081ff06",
        X"57558a76",
        X"27e2388b",
        X"19337f88",
        X"05349f19",
        X"339e1a33",
        X"71982b71",
        X"902b079d",
        X"1c337088",
        X"2b72079c",
        X"1e337107",
        X"640c5299",
        X"1d33981e",
        X"3371882b",
        X"07535153",
        X"57595674",
        X"7f840523",
        X"97193396",
        X"1a337188",
        X"2b075656",
        X"747f8605",
        X"23807734",
        X"7d51ebf0",
        X"3f83e080",
        X"08833270",
        X"30707207",
        X"9f2c83e0",
        X"80080652",
        X"5656961f",
        X"3355748a",
        X"38891f52",
        X"961f518d",
        X"9f3f7583",
        X"e0800c9e",
        X"3d0d04f4",
        X"3d0d7e8f",
        X"3dec1156",
        X"56589053",
        X"f0155277",
        X"51e0d23f",
        X"83e08008",
        X"80d63878",
        X"902e0981",
        X"0680cd38",
        X"02ab0533",
        X"80ece00b",
        X"80ece033",
        X"5758568c",
        X"3974762e",
        X"8a388417",
        X"70335657",
        X"74f33876",
        X"33705755",
        X"74802eac",
        X"38821722",
        X"708a2b90",
        X"3dec0556",
        X"70555656",
        X"96800a52",
        X"7751e081",
        X"3f83e080",
        X"08863878",
        X"752e8538",
        X"80568539",
        X"81173356",
        X"7583e080",
        X"0c8e3d0d",
        X"04fc3d0d",
        X"76705255",
        X"8ca63f83",
        X"e0800815",
        X"ff055473",
        X"752e8e38",
        X"73335372",
        X"ae2e8638",
        X"ff1454ef",
        X"39775281",
        X"14518bbe",
        X"3f83e080",
        X"08307083",
        X"e0800807",
        X"802583e0",
        X"800c5386",
        X"3d0d04fc",
        X"3d0d7670",
        X"5255e6ee",
        X"3f83e080",
        X"08548153",
        X"83e08008",
        X"80c13874",
        X"51e6b13f",
        X"83e08008",
        X"80ead053",
        X"83e08008",
        X"5253ff91",
        X"3f83e080",
        X"08a13880",
        X"ead45272",
        X"51ff823f",
        X"83e08008",
        X"923880ea",
        X"d8527251",
        X"fef33f83",
        X"e0800880",
        X"2e833881",
        X"54735372",
        X"83e0800c",
        X"863d0d04",
        X"fc3d0d76",
        X"705255e6",
        X"8d3f83e0",
        X"80085481",
        X"5383e080",
        X"0880d138",
        X"7451e5d0",
        X"3f83e080",
        X"0880ead0",
        X"5383e080",
        X"085253fe",
        X"b03f83e0",
        X"8008b138",
        X"80ead452",
        X"7251fea1",
        X"3f83e080",
        X"08a23880",
        X"ead85272",
        X"51fe923f",
        X"83e08008",
        X"933883e3",
        X"98085272",
        X"51fe823f",
        X"83e08008",
        X"802e8338",
        X"81547353",
        X"7283e080",
        X"0c863d0d",
        X"04fd3d0d",
        X"75705254",
        X"e59c3f81",
        X"5383e080",
        X"08983873",
        X"51e4e53f",
        X"83e38808",
        X"5283e080",
        X"0851fdc9",
        X"3f83e080",
        X"08537283",
        X"e0800c85",
        X"3d0d04df",
        X"3d0da43d",
        X"0870525e",
        X"db833f83",
        X"e0800833",
        X"953d5654",
        X"73963880",
        X"ede85274",
        X"5189ad3f",
        X"9a397d52",
        X"7851de8b",
        X"3f84ca39",
        X"7d51dae9",
        X"3f83e080",
        X"08527451",
        X"da993f80",
        X"43804280",
        X"41804083",
        X"e3900852",
        X"943d7052",
        X"5de0f33f",
        X"83e08008",
        X"59800b83",
        X"e0800855",
        X"5b83e080",
        X"087b2e94",
        X"38811b74",
        X"525be3f5",
        X"3f83e080",
        X"085483e0",
        X"8008ee38",
        X"805aff5f",
        X"7909709f",
        X"2c7b065b",
        X"547a7a24",
        X"8438ff1b",
        X"5af61a70",
        X"09709f2c",
        X"72067bff",
        X"125a5a52",
        X"55558075",
        X"25953876",
        X"51e3ba3f",
        X"83e08008",
        X"76ff1858",
        X"55577380",
        X"24ed3874",
        X"7f2e8638",
        X"a1e43f74",
        X"5f78ff1b",
        X"70585d58",
        X"807a2595",
        X"387751e3",
        X"903f83e0",
        X"800876ff",
        X"18585558",
        X"738024ed",
        X"38800b83",
        X"e7c00c80",
        X"0b83e7ec",
        X"0c80eadc",
        X"518dac3f",
        X"81800b83",
        X"e7ec0c80",
        X"eae4518d",
        X"9e3fa80b",
        X"83e7c00c",
        X"76802e80",
        X"e43883e7",
        X"c0087779",
        X"32703070",
        X"72078025",
        X"70872b83",
        X"e7ec0c51",
        X"56785356",
        X"56e2c73f",
        X"83e08008",
        X"802e8838",
        X"80eaec51",
        X"8ce53f76",
        X"51e2893f",
        X"83e08008",
        X"5280ec88",
        X"518cd43f",
        X"7651e291",
        X"3f83e080",
        X"0883e7c0",
        X"08555775",
        X"74258638",
        X"a81656f7",
        X"397583e7",
        X"c00c86f0",
        X"7624ff98",
        X"3887980b",
        X"83e7c00c",
        X"77802eb1",
        X"387751e1",
        X"c73f83e0",
        X"80087852",
        X"55e1e73f",
        X"80eaf454",
        X"83e08008",
        X"8d388739",
        X"80763481",
        X"ea3980ea",
        X"90547453",
        X"735280ea",
        X"f8518bf3",
        X"3f805480",
        X"eb80518b",
        X"ea3f8114",
        X"5473a82e",
        X"098106ef",
        X"38868da0",
        X"519dd83f",
        X"8052903d",
        X"705258b2",
        X"e73f8352",
        X"7751b2e0",
        X"3f6281ab",
        X"3861802e",
        X"8197387b",
        X"5473ff2e",
        X"96387880",
        X"2e818638",
        X"7851e0ed",
        X"3f83e080",
        X"08ff1555",
        X"59e73978",
        X"802e80f1",
        X"387851e0",
        X"e93f83e0",
        X"8008802e",
        X"fc903878",
        X"51e0b13f",
        X"83e08008",
        X"5280eacc",
        X"5184823f",
        X"83e08008",
        X"bb387c51",
        X"85ba3f83",
        X"e08008ff",
        X"0555800b",
        X"83e08008",
        X"2580c838",
        X"a33d7505",
        X"c4057058",
        X"567633ff",
        X"18585473",
        X"af2efec4",
        X"3874ff16",
        X"ff185856",
        X"54738024",
        X"e838a439",
        X"7851dfda",
        X"3f83e080",
        X"08527c51",
        X"84da3f93",
        X"3981549e",
        X"397f1060",
        X"8829057a",
        X"0561055a",
        X"fbf63962",
        X"802efbb7",
        X"38805277",
        X"51b1a53f",
        X"80547383",
        X"e0800ca3",
        X"3d0d0480",
        X"3d0d9088",
        X"b8337081",
        X"ff067084",
        X"2a813270",
        X"81065151",
        X"51517080",
        X"2e8d38a8",
        X"0b9088b8",
        X"34b80b90",
        X"88b83470",
        X"83e0800c",
        X"823d0d04",
        X"803d0d90",
        X"88b83370",
        X"81ff0670",
        X"852a8132",
        X"70810651",
        X"51515170",
        X"802e8d38",
        X"980b9088",
        X"b834b80b",
        X"9088b834",
        X"7083e080",
        X"0c823d0d",
        X"04930b90",
        X"88bc34ff",
        X"0b9088a8",
        X"3404ff3d",
        X"0d028f05",
        X"3352800b",
        X"9088bc34",
        X"8a519aff",
        X"3fdf3f80",
        X"f80b9088",
        X"a034800b",
        X"90888834",
        X"fa125271",
        X"90888034",
        X"800b9088",
        X"98347190",
        X"88903490",
        X"88b85280",
        X"7234b872",
        X"34833d0d",
        X"04803d0d",
        X"028b0533",
        X"51709088",
        X"b434febf",
        X"3f83e080",
        X"08802ef6",
        X"38823d0d",
        X"04803d0d",
        X"8439a8ab",
        X"3ffed93f",
        X"83e08008",
        X"802ef338",
        X"9088b433",
        X"7081ff06",
        X"83e0800c",
        X"51823d0d",
        X"04803d0d",
        X"a30b9088",
        X"bc34ff0b",
        X"9088a834",
        X"9088b851",
        X"a87134b8",
        X"7134823d",
        X"0d04803d",
        X"0d9088bc",
        X"3370982b",
        X"70802583",
        X"e0800c51",
        X"51823d0d",
        X"04803d0d",
        X"9088b833",
        X"7081ff06",
        X"70832a81",
        X"32708106",
        X"51515151",
        X"70802ee8",
        X"38b00b90",
        X"88b834b8",
        X"0b9088b8",
        X"34823d0d",
        X"04803d0d",
        X"9080ac08",
        X"810683e0",
        X"800c823d",
        X"0d04fd3d",
        X"0d757754",
        X"54807325",
        X"94387370",
        X"81055533",
        X"5280eb84",
        X"5187843f",
        X"ff1353e9",
        X"39853d0d",
        X"04fd3d0d",
        X"75775354",
        X"73335170",
        X"89387133",
        X"5170802e",
        X"a1387333",
        X"72335253",
        X"72712785",
        X"38ff5194",
        X"39707327",
        X"85388151",
        X"8b398114",
        X"81135354",
        X"d3398051",
        X"7083e080",
        X"0c853d0d",
        X"04fd3d0d",
        X"75775454",
        X"72337081",
        X"ff065252",
        X"70802ea3",
        X"387181ff",
        X"068114ff",
        X"bf125354",
        X"52709926",
        X"8938a012",
        X"7081ff06",
        X"53517174",
        X"70810556",
        X"34d23980",
        X"7434853d",
        X"0d04ffbd",
        X"3d0d80c6",
        X"3d0852a5",
        X"3d705254",
        X"ffb33f80",
        X"c73d0852",
        X"853d7052",
        X"53ffa63f",
        X"72527351",
        X"fedf3f80",
        X"c53d0d04",
        X"fe3d0d74",
        X"76535371",
        X"70810553",
        X"33517073",
        X"70810555",
        X"3470f038",
        X"843d0d04",
        X"fe3d0d74",
        X"52807233",
        X"52537073",
        X"2e8d3881",
        X"12811471",
        X"33535452",
        X"70f53872",
        X"83e0800c",
        X"843d0d04",
        X"f63d0d7c",
        X"7e60625a",
        X"5d5b5680",
        X"59815585",
        X"39747a29",
        X"55745275",
        X"51ad833f",
        X"83e08008",
        X"7a27ee38",
        X"74802e80",
        X"dd387452",
        X"7551acee",
        X"3f83e080",
        X"08755376",
        X"5254acf2",
        X"3f83e080",
        X"087a5375",
        X"5256acd6",
        X"3f83e080",
        X"08793070",
        X"7b079f2a",
        X"70778024",
        X"07515154",
        X"55728738",
        X"83e08008",
        X"c5387681",
        X"18b01655",
        X"58588974",
        X"258b38b7",
        X"14537a85",
        X"3880d714",
        X"53727834",
        X"811959ff",
        X"9f398077",
        X"348c3d0d",
        X"04f73d0d",
        X"7b7d7f62",
        X"029005bb",
        X"05335759",
        X"565a5ab0",
        X"58728338",
        X"a0587570",
        X"70810552",
        X"33715954",
        X"55903980",
        X"74258e38",
        X"ff147770",
        X"81055933",
        X"545472ef",
        X"3873ff15",
        X"55538073",
        X"25893877",
        X"52795178",
        X"2def3975",
        X"33755753",
        X"72802e90",
        X"38725279",
        X"51782d75",
        X"70810557",
        X"3353ed39",
        X"8b3d0d04",
        X"ee3d0d64",
        X"66696970",
        X"70810552",
        X"335b4a5c",
        X"5e5e7680",
        X"2e82f938",
        X"76a52e09",
        X"810682e0",
        X"38807041",
        X"67707081",
        X"05523371",
        X"4a59575f",
        X"76b02e09",
        X"81068c38",
        X"75708105",
        X"57337648",
        X"57815fd0",
        X"17567589",
        X"2680da38",
        X"76675c59",
        X"805c9339",
        X"778a2480",
        X"c3387b8a",
        X"29187b70",
        X"81055d33",
        X"5a5cd019",
        X"7081ff06",
        X"58588977",
        X"27a438ff",
        X"9f197081",
        X"ff06ffa9",
        X"1b5a5156",
        X"85762792",
        X"38ffbf19",
        X"7081ff06",
        X"51567585",
        X"268a38c9",
        X"19587780",
        X"25ffb938",
        X"7a477b40",
        X"7881ff06",
        X"577680e4",
        X"2e80e538",
        X"7680e424",
        X"a7387680",
        X"d82e8186",
        X"387680d8",
        X"24903876",
        X"802e81cc",
        X"3876a52e",
        X"81b63881",
        X"b9397680",
        X"e32e818c",
        X"3881af39",
        X"7680f52e",
        X"9b387680",
        X"f5248b38",
        X"7680f32e",
        X"81813881",
        X"99397680",
        X"f82e80ca",
        X"38818f39",
        X"913d7055",
        X"5780538a",
        X"5279841b",
        X"7108535b",
        X"56fc813f",
        X"7655ab39",
        X"79841b71",
        X"08943d70",
        X"5b5b525b",
        X"56758025",
        X"8c387530",
        X"56ad7834",
        X"0280c105",
        X"57765480",
        X"538a5275",
        X"51fbd53f",
        X"77557e54",
        X"b839913d",
        X"70557780",
        X"d8327030",
        X"70802556",
        X"51585690",
        X"5279841b",
        X"7108535b",
        X"57fbb13f",
        X"7555db39",
        X"79841b83",
        X"1233545b",
        X"56983979",
        X"841b7108",
        X"575b5680",
        X"547f537c",
        X"527d51fc",
        X"9c3f8739",
        X"76527d51",
        X"7c2d6670",
        X"33588105",
        X"47fd8339",
        X"943d0d04",
        X"7283e094",
        X"0c7183e0",
        X"980c04fb",
        X"3d0d883d",
        X"70708405",
        X"52085754",
        X"755383e0",
        X"94085283",
        X"e0980851",
        X"fcc63f87",
        X"3d0d04ff",
        X"3d0d7370",
        X"08535102",
        X"93053372",
        X"34700881",
        X"05710c83",
        X"3d0d04fc",
        X"3d0d873d",
        X"88115578",
        X"54becf53",
        X"51fc993f",
        X"8052873d",
        X"51d13f86",
        X"3d0d04fc",
        X"3d0d7655",
        X"7483e39c",
        X"082eaf38",
        X"80537451",
        X"87c63f83",
        X"e0800881",
        X"ff06ff14",
        X"7081ff06",
        X"7230709f",
        X"2a515255",
        X"53547280",
        X"2e843871",
        X"dd3873fe",
        X"387483e3",
        X"9c0c863d",
        X"0d04ff3d",
        X"0dff0b83",
        X"e39c0c84",
        X"a53f8151",
        X"878a3f83",
        X"e0800881",
        X"ff065271",
        X"ee3881d3",
        X"3f7183e0",
        X"800c833d",
        X"0d04fc3d",
        X"0d760284",
        X"05a20522",
        X"028805a6",
        X"05227a54",
        X"555555ff",
        X"823f7280",
        X"2ea03883",
        X"e3b01433",
        X"75708105",
        X"57348114",
        X"7083ffff",
        X"06ff1570",
        X"83ffff06",
        X"56525552",
        X"dd39800b",
        X"83e0800c",
        X"863d0d04",
        X"fc3d0d76",
        X"787a1156",
        X"53558053",
        X"71742e93",
        X"38741351",
        X"703383e3",
        X"b0133481",
        X"12811454",
        X"52ea3980",
        X"0b83e080",
        X"0c863d0d",
        X"04fd3d0d",
        X"905483e3",
        X"9c085186",
        X"f93f83e0",
        X"800881ff",
        X"06ff1571",
        X"30713070",
        X"73079f2a",
        X"729f2a06",
        X"52555255",
        X"5372db38",
        X"853d0d04",
        X"803d0d83",
        X"e3a80810",
        X"83e3a008",
        X"079080a8",
        X"0c823d0d",
        X"04800b83",
        X"e3a80ce4",
        X"3f04810b",
        X"83e3a80c",
        X"db3f04ed",
        X"3f047183",
        X"e3a40c04",
        X"803d0d80",
        X"51f43f81",
        X"0b83e3a8",
        X"0c810b83",
        X"e3a00cff",
        X"bb3f823d",
        X"0d04803d",
        X"0d723070",
        X"74078025",
        X"83e3a00c",
        X"51ffa53f",
        X"823d0d04",
        X"803d0d02",
        X"8b053390",
        X"80a40c90",
        X"80a80870",
        X"81065151",
        X"70f53890",
        X"80a40870",
        X"81ff0683",
        X"e0800c51",
        X"823d0d04",
        X"803d0d81",
        X"ff51d13f",
        X"83e08008",
        X"81ff0683",
        X"e0800c82",
        X"3d0d0480",
        X"3d0d7390",
        X"2b730790",
        X"80b40c82",
        X"3d0d0404",
        X"fb3d0d78",
        X"0284059f",
        X"05337098",
        X"2b555755",
        X"7280259b",
        X"387580ff",
        X"06568052",
        X"80f751e0",
        X"3f83e080",
        X"0881ff06",
        X"54738126",
        X"80ff3880",
        X"51fee73f",
        X"ffa23f81",
        X"51fedf3f",
        X"ff9a3f75",
        X"51feed3f",
        X"74982a51",
        X"fee63f74",
        X"902a7081",
        X"ff065253",
        X"feda3f74",
        X"882a7081",
        X"ff065253",
        X"fece3f74",
        X"81ff0651",
        X"fec63f81",
        X"557580c0",
        X"2e098106",
        X"86388195",
        X"558d3975",
        X"80c82e09",
        X"81068438",
        X"81875574",
        X"51fea53f",
        X"8a55fec8",
        X"3f83e080",
        X"0881ff06",
        X"70982b54",
        X"54728025",
        X"8c38ff15",
        X"7081ff06",
        X"565374e2",
        X"387383e0",
        X"800c873d",
        X"0d04fa3d",
        X"0dfdc53f",
        X"8051fdda",
        X"3f8a54fe",
        X"933fff14",
        X"7081ff06",
        X"555373f3",
        X"38737453",
        X"5580c051",
        X"fea63f83",
        X"e0800881",
        X"ff065473",
        X"812e0981",
        X"0682a438",
        X"83aa5280",
        X"c851fe8c",
        X"3f83e080",
        X"0881ff06",
        X"5372812e",
        X"09810681",
        X"ad387454",
        X"883d7405",
        X"fc0553fd",
        X"c73f83e0",
        X"80087334",
        X"81147081",
        X"ff065553",
        X"837427e4",
        X"38029a05",
        X"33537281",
        X"2e098106",
        X"81dd3802",
        X"9b053353",
        X"80ce9054",
        X"7281aa2e",
        X"8d3881cb",
        X"3980e451",
        X"8ba93fff",
        X"14547380",
        X"2e81bc38",
        X"820a5281",
        X"e951fda4",
        X"3f83e080",
        X"0881ff06",
        X"5372de38",
        X"725280fa",
        X"51fd913f",
        X"83e08008",
        X"81ff0653",
        X"72819438",
        X"7254883d",
        X"7405fc05",
        X"53fcd13f",
        X"83e08008",
        X"73348114",
        X"7081ff06",
        X"55538374",
        X"27e43887",
        X"3d337086",
        X"2a708106",
        X"5154568c",
        X"557280e3",
        X"38845580",
        X"de397452",
        X"81e951fc",
        X"c73f83e0",
        X"800881ff",
        X"06538255",
        X"81e95681",
        X"73278638",
        X"735580c1",
        X"5680ce90",
        X"548a3980",
        X"e4518a97",
        X"3fff1454",
        X"73802ea9",
        X"38805275",
        X"51fc953f",
        X"83e08008",
        X"81ff0653",
        X"72e13884",
        X"805280d0",
        X"51fc813f",
        X"83e08008",
        X"81ff0653",
        X"72802e83",
        X"38805574",
        X"83e3ac34",
        X"8051fb82",
        X"3ffbbd3f",
        X"883d0d04",
        X"fb3d0d77",
        X"54800b83",
        X"e3ac3370",
        X"832a7081",
        X"06515557",
        X"5572752e",
        X"09810685",
        X"3873892b",
        X"54735280",
        X"d151fbb8",
        X"3f83e080",
        X"0881ff06",
        X"5372bd38",
        X"82b8c054",
        X"fafe3f83",
        X"e0800881",
        X"ff065372",
        X"81ff2e09",
        X"81068938",
        X"ff145473",
        X"e7389f39",
        X"7281fe2e",
        X"09810696",
        X"3883e7b0",
        X"5283e3b0",
        X"51fae83f",
        X"face3ffa",
        X"cb3f8339",
        X"81558051",
        X"fa843ffa",
        X"bf3f7481",
        X"ff0683e0",
        X"800c873d",
        X"0d04fb3d",
        X"0d7783e3",
        X"b0565481",
        X"51f9e73f",
        X"83e3ac33",
        X"70832a70",
        X"81065154",
        X"56728538",
        X"73892b54",
        X"735280d8",
        X"51fab13f",
        X"83e08008",
        X"81ff0653",
        X"7280e438",
        X"81ff51f9",
        X"cf3f81fe",
        X"51f9c93f",
        X"84805374",
        X"70810556",
        X"3351f9bc",
        X"3fff1370",
        X"83ffff06",
        X"515372eb",
        X"387251f9",
        X"ab3f7251",
        X"f9a63ff9",
        X"cb3f83e0",
        X"80089f06",
        X"53a78854",
        X"72852e8c",
        X"38993980",
        X"e45187cf",
        X"3fff1454",
        X"f9ae3f83",
        X"e0800881",
        X"ff2e8438",
        X"73e93880",
        X"51f8df3f",
        X"f99a3f80",
        X"0b83e080",
        X"0c873d0d",
        X"047183e7",
        X"b40c8880",
        X"800b83e7",
        X"b00c8480",
        X"800b83e7",
        X"b80c04f1",
        X"3d0d8380",
        X"805683e7",
        X"b4081683",
        X"e7b00817",
        X"56547433",
        X"743483e7",
        X"b8081654",
        X"80743481",
        X"16567583",
        X"80a02e09",
        X"8106db38",
        X"83d08056",
        X"83e7b408",
        X"1683e7b0",
        X"08175654",
        X"74337434",
        X"83e7b808",
        X"16548074",
        X"34811656",
        X"7583d090",
        X"2e098106",
        X"db3883a8",
        X"805683e7",
        X"b4081683",
        X"e7b00817",
        X"56547433",
        X"743483e7",
        X"b8081654",
        X"80743481",
        X"16567583",
        X"a8902e09",
        X"8106db38",
        X"805683e7",
        X"b4081683",
        X"e7b80817",
        X"55557333",
        X"75348116",
        X"56758180",
        X"802e0981",
        X"06e43887",
        X"f53f883d",
        X"54a25380",
        X"ea945273",
        X"519e873f",
        X"80558c80",
        X"74585683",
        X"e7b80816",
        X"54767081",
        X"05583374",
        X"34811681",
        X"16565674",
        X"a22e0981",
        X"06e53886",
        X"0b87a883",
        X"34800b87",
        X"a8823480",
        X"0b87809a",
        X"34af0b87",
        X"809634bf",
        X"0b878097",
        X"34800b87",
        X"8098349f",
        X"0b878099",
        X"34800b87",
        X"809b34f8",
        X"0b87a889",
        X"347487a8",
        X"8034820b",
        X"87d08f34",
        X"820b87a8",
        X"8134840b",
        X"87809f34",
        X"ff0b87d0",
        X"8b34913d",
        X"0d04fe3d",
        X"0d805383",
        X"e7b80813",
        X"83e7b408",
        X"14525270",
        X"33723481",
        X"13537281",
        X"80802e09",
        X"8106e438",
        X"83808053",
        X"83e7b808",
        X"1383e7b4",
        X"08145252",
        X"70337234",
        X"81135372",
        X"8380a02e",
        X"098106e4",
        X"3883d080",
        X"5383e7b8",
        X"081383e7",
        X"b4081452",
        X"52703372",
        X"34811353",
        X"7283d090",
        X"2e098106",
        X"e43883a8",
        X"805383e7",
        X"b8081383",
        X"e7b40814",
        X"52527033",
        X"72348113",
        X"537283a8",
        X"902e0981",
        X"06e43884",
        X"3d0d0480",
        X"3d0d9080",
        X"90088106",
        X"83e0800c",
        X"823d0d04",
        X"ff3d0d90",
        X"80907008",
        X"70fe0676",
        X"07720c52",
        X"52833d0d",
        X"04803d0d",
        X"90809008",
        X"70812c81",
        X"0683e080",
        X"0c51823d",
        X"0d04ff3d",
        X"0d908090",
        X"700870fd",
        X"06761007",
        X"720c5252",
        X"833d0d04",
        X"803d0d90",
        X"80900870",
        X"822cbf06",
        X"83e0800c",
        X"51823d0d",
        X"04ff3d0d",
        X"90809070",
        X"0870fe83",
        X"0676822b",
        X"07720c52",
        X"52833d0d",
        X"04803d0d",
        X"90809008",
        X"70882c87",
        X"0683e080",
        X"0c51823d",
        X"0d04ff3d",
        X"0d908090",
        X"700870f1",
        X"ff067688",
        X"2b07720c",
        X"5252833d",
        X"0d04803d",
        X"0d908090",
        X"0870912c",
        X"bf0683e0",
        X"800c5182",
        X"3d0d04ff",
        X"3d0d9080",
        X"90700870",
        X"fc87ffff",
        X"0676912b",
        X"07720c52",
        X"52833d0d",
        X"04803d0d",
        X"90809008",
        X"70992c81",
        X"0683e080",
        X"0c51823d",
        X"0d04ff3d",
        X"0d908090",
        X"700870ff",
        X"bf0a0676",
        X"992b0772",
        X"0c525283",
        X"3d0d0480",
        X"3d0d9080",
        X"9008709a",
        X"2c810683",
        X"e0800c51",
        X"823d0d04",
        X"ff3d0d90",
        X"80907008",
        X"70df0a06",
        X"769a2b07",
        X"720c5252",
        X"833d0d04",
        X"803d0d90",
        X"80900870",
        X"9b2c8106",
        X"83e0800c",
        X"51823d0d",
        X"04ff3d0d",
        X"90809070",
        X"0870ef0a",
        X"06769b2b",
        X"07720c52",
        X"52833d0d",
        X"04803d0d",
        X"90808008",
        X"70882c81",
        X"0683e080",
        X"0c51823d",
        X"0d04803d",
        X"0d908080",
        X"0870892c",
        X"810683e0",
        X"800c5182",
        X"3d0d0480",
        X"3d0d9080",
        X"8008708a",
        X"2c810683",
        X"e0800c51",
        X"823d0d04",
        X"803d0d90",
        X"80800870",
        X"8b2c8106",
        X"83e0800c",
        X"51823d0d",
        X"04803d0d",
        X"90808008",
        X"70922c81",
        X"0683e080",
        X"0c51823d",
        X"0d04803d",
        X"0d908080",
        X"08708c2c",
        X"bf0683e0",
        X"800c5182",
        X"3d0d04fe",
        X"3d0d7481",
        X"e629872a",
        X"9080a00c",
        X"843d0d04",
        X"fe3d0d75",
        X"75ff1953",
        X"535370ff",
        X"2e8d3872",
        X"72708105",
        X"5434ff11",
        X"51f03984",
        X"3d0d04fe",
        X"3d0d7575",
        X"ff195353",
        X"5370ff2e",
        X"8d387272",
        X"70840554",
        X"0cff1151",
        X"f039843d",
        X"0d04fe3d",
        X"0d818080",
        X"53805288",
        X"800a51ff",
        X"b33fa080",
        X"53805282",
        X"800a51c7",
        X"3f843d0d",
        X"04803d0d",
        X"8151fbbc",
        X"3f72802e",
        X"90388051",
        X"fd903fce",
        X"3f80edd4",
        X"3351fd86",
        X"3f8151fb",
        X"cd3f8051",
        X"fbc83f80",
        X"51fb993f",
        X"823d0d04",
        X"fd3d0d75",
        X"52805480",
        X"ff722588",
        X"38810bff",
        X"80135354",
        X"ffbf1251",
        X"70992686",
        X"38e01252",
        X"b039ff9f",
        X"12519971",
        X"27a738d0",
        X"12e01354",
        X"51708926",
        X"85387252",
        X"9839728f",
        X"26853872",
        X"528f3971",
        X"ba2e0981",
        X"0685389a",
        X"52833980",
        X"5273802e",
        X"85388180",
        X"12527181",
        X"ff0683e0",
        X"800c853d",
        X"0d04803d",
        X"0d84d8c0",
        X"51807170",
        X"81055334",
        X"7084e0c0",
        X"2e098106",
        X"f038823d",
        X"0d04fe3d",
        X"0d029705",
        X"3351fef4",
        X"3f83e080",
        X"0881ff06",
        X"83e7c008",
        X"54528073",
        X"249b3883",
        X"e7e80813",
        X"7283e7ec",
        X"08075353",
        X"71733483",
        X"e7c00881",
        X"0583e7c0",
        X"0c843d0d",
        X"04fa3d0d",
        X"82800a1b",
        X"55805788",
        X"3dfc0554",
        X"79537452",
        X"7851ffb9",
        X"8c3f883d",
        X"0d04fe3d",
        X"0d83e7d8",
        X"08527451",
        X"ffbfef3f",
        X"83e08008",
        X"8c387653",
        X"755283e7",
        X"d80851c5",
        X"3f843d0d",
        X"04fe3d0d",
        X"83e7d808",
        X"53755274",
        X"51ffbaad",
        X"3f83e080",
        X"088d3877",
        X"53765283",
        X"e7d80851",
        X"ff9f3f84",
        X"3d0d04fd",
        X"3d0d83e7",
        X"d80851ff",
        X"b9a03f83",
        X"e0800890",
        X"802e0981",
        X"06ad3880",
        X"5483c180",
        X"805383e0",
        X"80085283",
        X"e7d80851",
        X"feef3f87",
        X"c1808014",
        X"3387c190",
        X"80153481",
        X"14547390",
        X"802e0981",
        X"06e93885",
        X"3d0d04fc",
        X"3d0d7654",
        X"73902e80",
        X"ff387390",
        X"248e3873",
        X"842e9838",
        X"73862ea6",
        X"3882b939",
        X"73932e81",
        X"95387394",
        X"2e81cf38",
        X"82aa3981",
        X"80805382",
        X"80805283",
        X"e7d40851",
        X"fe973f82",
        X"b5398054",
        X"81808053",
        X"80c08052",
        X"83e7d408",
        X"51fe823f",
        X"82808053",
        X"80c08052",
        X"83e7d408",
        X"51fdf23f",
        X"84818080",
        X"14338481",
        X"c0801534",
        X"84828080",
        X"14338482",
        X"c0801534",
        X"81145473",
        X"80c0802e",
        X"098106dc",
        X"3881eb39",
        X"82808053",
        X"81808052",
        X"83e7d408",
        X"51fdba3f",
        X"80548482",
        X"80801433",
        X"84818080",
        X"15348114",
        X"54738180",
        X"802e0981",
        X"06e83881",
        X"bd398180",
        X"805380c0",
        X"805283e7",
        X"d40851fd",
        X"8c3f8055",
        X"84818080",
        X"15547333",
        X"8481c080",
        X"16347333",
        X"84828080",
        X"16347333",
        X"8482c080",
        X"16348115",
        X"557480c0",
        X"802e0981",
        X"06d63880",
        X"fd398180",
        X"8053a080",
        X"5283e7d4",
        X"0851fccd",
        X"3f805584",
        X"81808015",
        X"54733384",
        X"81a08016",
        X"34733384",
        X"81c08016",
        X"34733384",
        X"81e08016",
        X"34733384",
        X"82808016",
        X"34733384",
        X"82a08016",
        X"34733384",
        X"82c08016",
        X"34733384",
        X"82e08016",
        X"34811555",
        X"74a0802e",
        X"098106ff",
        X"b6389f39",
        X"fba43f80",
        X"0b83e7c0",
        X"0c800b83",
        X"e7ec0c80",
        X"eb8c51e7",
        X"8e3f81b7",
        X"8dc051f9",
        X"863f863d",
        X"0d04fc3d",
        X"0d767052",
        X"55ffbcca",
        X"3f83e080",
        X"08548153",
        X"83e08008",
        X"80c23874",
        X"51ffbc8c",
        X"3f83e080",
        X"0880eba8",
        X"5383e080",
        X"085253d4",
        X"ec3f83e0",
        X"8008a138",
        X"80ebac52",
        X"7251d4dd",
        X"3f83e080",
        X"08923880",
        X"ebb05272",
        X"51d4ce3f",
        X"83e08008",
        X"802e8338",
        X"81547353",
        X"7283e080",
        X"0c863d0d",
        X"04f13d0d",
        X"80d7ae0b",
        X"83e3900c",
        X"83e7d408",
        X"51d6ec3f",
        X"83e08008",
        X"5583e080",
        X"08802e81",
        X"ea3883e7",
        X"d40851ff",
        X"b1e33fff",
        X"0b80ebac",
        X"5383e080",
        X"085256d4",
        X"803f83e0",
        X"8008802e",
        X"9f388058",
        X"913ddc11",
        X"55559053",
        X"f0155283",
        X"e7d40851",
        X"ffb3c63f",
        X"02b70533",
        X"5681a539",
        X"83e7d408",
        X"51ffb4a2",
        X"3f83e080",
        X"085783e0",
        X"80088280",
        X"802e0981",
        X"06833884",
        X"5683e080",
        X"08818080",
        X"2e098106",
        X"80e13880",
        X"5c805b80",
        X"5a8059f9",
        X"8d3f800b",
        X"83e7c00c",
        X"800b83e7",
        X"ec0c80eb",
        X"b451e4f7",
        X"3f80d00b",
        X"83e7c00c",
        X"80ebc451",
        X"e4e93f80",
        X"f80b83e7",
        X"c00c80eb",
        X"d851e4db",
        X"3f758025",
        X"a2388052",
        X"893d7052",
        X"558be53f",
        X"83527451",
        X"8bde3f78",
        X"55748025",
        X"83389056",
        X"807525dd",
        X"38865676",
        X"80c0802e",
        X"09810685",
        X"3893568c",
        X"3976a080",
        X"2e098106",
        X"83389456",
        X"7551fa9f",
        X"3f815574",
        X"83e0800c",
        X"913d0d04",
        X"f73d0d80",
        X"5a805980",
        X"58805780",
        X"705656f7",
        X"fd3f800b",
        X"83e7c00c",
        X"800b83e7",
        X"ec0c80eb",
        X"ec51e3e7",
        X"3f81800b",
        X"83e7ec0c",
        X"80ebf051",
        X"e3d93f80",
        X"d00b83e7",
        X"c00c7430",
        X"70760780",
        X"2570872b",
        X"83e7ec0c",
        X"5153f2b0",
        X"3f83e080",
        X"085280eb",
        X"f851e3b3",
        X"3f80f80b",
        X"83e7c00c",
        X"74813270",
        X"30707207",
        X"80257087",
        X"2b83e7ec",
        X"0c515483",
        X"e7d80852",
        X"54ffaefd",
        X"3f83e080",
        X"085280ec",
        X"8451e383",
        X"3f81a00b",
        X"83e7c00c",
        X"74823270",
        X"30707207",
        X"80257087",
        X"2b83e7ec",
        X"0c515483",
        X"e7d40852",
        X"54ffaecd",
        X"3f80ec8c",
        X"5383e080",
        X"08802e8f",
        X"3883e7d4",
        X"0851ffae",
        X"b83f83e0",
        X"80085372",
        X"5280ec94",
        X"51e2bc3f",
        X"81f00b83",
        X"e7c00c74",
        X"83327030",
        X"70720780",
        X"2570872b",
        X"83e7ec0c",
        X"515454f2",
        X"c63f80ec",
        X"9c5383e0",
        X"80088538",
        X"80eca053",
        X"725280ec",
        X"a851e287",
        X"3f82c00b",
        X"83e7c00c",
        X"74843270",
        X"30707207",
        X"80257087",
        X"2b83e7ec",
        X"0c515580",
        X"ecbc5253",
        X"e1e53f86",
        X"8da051f3",
        X"de3f8052",
        X"873d7052",
        X"5388ed3f",
        X"83527251",
        X"88e63f79",
        X"537281bc",
        X"38771555",
        X"74802585",
        X"38845590",
        X"39847525",
        X"85387255",
        X"87397484",
        X"26819b38",
        X"74842980",
        X"eab80553",
        X"720804f0",
        X"8f3f83e0",
        X"80087755",
        X"5373812e",
        X"09810689",
        X"3883e080",
        X"08105390",
        X"3973ff2e",
        X"09810688",
        X"3883e080",
        X"08812c53",
        X"90732585",
        X"38905388",
        X"39728024",
        X"83388153",
        X"7251efe9",
        X"3f80cf39",
        X"76873878",
        X"802e80c6",
        X"3883e38c",
        X"0883e388",
        X"0caedd0b",
        X"83e3900c",
        X"83e7d808",
        X"51d1a03f",
        X"f5fd3faa",
        X"39768638",
        X"78802ea2",
        X"38fa923f",
        X"83e08008",
        X"53a03976",
        X"802e9338",
        X"f0c93f83",
        X"e0800881",
        X"3251f0d4",
        X"3f843978",
        X"87387580",
        X"2efc9038",
        X"80537283",
        X"e0800c8b",
        X"3d0d04f9",
        X"3d0d8058",
        X"80578056",
        X"8055f0f5",
        X"3f83e080",
        X"08802e86",
        X"38805180",
        X"f839f0fa",
        X"3f83e080",
        X"0880ec38",
        X"f19a3f83",
        X"e0800880",
        X"2eb43881",
        X"51edfd3f",
        X"eab53f80",
        X"0b83e7c0",
        X"0cfbb53f",
        X"83e08008",
        X"53805289",
        X"3df00551",
        X"86ca3fff",
        X"0b83e7c0",
        X"0cecbf3f",
        X"72b53872",
        X"51edd13f",
        X"b339f0c7",
        X"3f83e080",
        X"08802ea8",
        X"388151ed",
        X"bf3fe9f7",
        X"3ff8ea3f",
        X"83e08008",
        X"53805289",
        X"3df00551",
        X"86923fec",
        X"8d3f7280",
        X"2e863881",
        X"51f1da3f",
        X"893d0d04",
        X"fe3d0d82",
        X"80805380",
        X"52818180",
        X"8051f0e8",
        X"3f80c080",
        X"53805284",
        X"81808051",
        X"f0f93f90",
        X"80805286",
        X"84808051",
        X"ffaed03f",
        X"83e08008",
        X"a43880ed",
        X"d851ffb3",
        X"933f83e7",
        X"d8085380",
        X"ecc45283",
        X"e0800851",
        X"ffadf23f",
        X"83e08008",
        X"8438f3d3",
        X"3f8151f0",
        X"fc3ffe8b",
        X"3ffc3983",
        X"e08c0802",
        X"83e08c0c",
        X"fb3d0d02",
        X"80ecd00b",
        X"83e38c0c",
        X"80ebb00b",
        X"83e3840c",
        X"80ebac0b",
        X"83e3980c",
        X"80ecd40b",
        X"83e3940c",
        X"83e08c08",
        X"fc050c80",
        X"0b83e7c4",
        X"0b83e08c",
        X"08f8050c",
        X"83e08c08",
        X"f4050cff",
        X"acc93f83",
        X"e0800886",
        X"05fc0683",
        X"e08c08f0",
        X"050c0283",
        X"e08c08f0",
        X"0508310d",
        X"833d7083",
        X"e08c08f8",
        X"05087084",
        X"0583e08c",
        X"08f8050c",
        X"0c51ffa9",
        X"8a3f83e0",
        X"8c08f405",
        X"08810583",
        X"e08c08f4",
        X"050c83e0",
        X"8c08f405",
        X"08892e09",
        X"8106ffab",
        X"38869480",
        X"8051e7b9",
        X"3fff0b83",
        X"e7c00c80",
        X"0b83e7ec",
        X"0c84d8c0",
        X"0b83e7e8",
        X"0c8151ea",
        X"fb3f8151",
        X"eba03f80",
        X"51eb9b3f",
        X"ebae3f83",
        X"e080088b",
        X"388151eb",
        X"b83f8251",
        X"ebe03f80",
        X"51ec883f",
        X"8051ecb2",
        X"3f80d2ce",
        X"528051dc",
        X"8f3ffdb0",
        X"3f83e08c",
        X"08fc0508",
        X"0d800b83",
        X"e0800c87",
        X"3d0d83e0",
        X"8c0c04fb",
        X"3d0d7754",
        X"80740c80",
        X"0b84150c",
        X"800b8815",
        X"0c800b8c",
        X"150cedd2",
        X"3f83e080",
        X"0887d088",
        X"337081ff",
        X"06515255",
        X"70a73887",
        X"d0803383",
        X"e7fc3487",
        X"d0813383",
        X"e7f83487",
        X"d0823383",
        X"e7f03487",
        X"d0833383",
        X"e7f434ff",
        X"0b87d08b",
        X"3487d089",
        X"3387d08f",
        X"3370822a",
        X"70810670",
        X"30707207",
        X"7009709f",
        X"2c77069e",
        X"06575151",
        X"55515153",
        X"53807398",
        X"06525270",
        X"882e0981",
        X"06833881",
        X"52709832",
        X"70307080",
        X"25747131",
        X"84180c51",
        X"51518073",
        X"86065252",
        X"70822e09",
        X"81068338",
        X"81527086",
        X"32703070",
        X"80257471",
        X"31770c51",
        X"515183e7",
        X"fc335181",
        X"aa712784",
        X"3881740c",
        X"83e7fc33",
        X"5170bb26",
        X"8438ff74",
        X"0c83e7f8",
        X"335181aa",
        X"71278638",
        X"810b8415",
        X"0c83e7f8",
        X"335170bb",
        X"268638ff",
        X"0b84150c",
        X"83e7f033",
        X"5181aa71",
        X"27843881",
        X"740c83e7",
        X"f0335170",
        X"bb268438",
        X"ff740c83",
        X"e7f43351",
        X"81aa7127",
        X"8638810b",
        X"84150c83",
        X"e7f43351",
        X"70bb2686",
        X"38ff0b84",
        X"150c8056",
        X"72942eaa",
        X"38878090",
        X"33878091",
        X"33878092",
        X"337081ff",
        X"06727406",
        X"06878093",
        X"33710681",
        X"06515253",
        X"53537176",
        X"2e098106",
        X"83388156",
        X"7588150c",
        X"74802eb0",
        X"3874812a",
        X"70810676",
        X"81063184",
        X"160c5174",
        X"832a7582",
        X"2a718106",
        X"71810631",
        X"760c5252",
        X"74842a81",
        X"0688150c",
        X"74852a81",
        X"068c150c",
        X"873d0d04",
        X"fe3d0d74",
        X"76545271",
        X"51fcdc3f",
        X"ea9a3f83",
        X"e0800880",
        X"2e893881",
        X"0b8c130c",
        X"80d03972",
        X"812ea738",
        X"8173268d",
        X"3872822e",
        X"ad387283",
        X"2ea138d3",
        X"397108cf",
        X"38841208",
        X"ca388812",
        X"08c5388c",
        X"1208c038",
        X"a5398812",
        X"08812e9e",
        X"38913988",
        X"1208812e",
        X"95387108",
        X"91388412",
        X"088c388c",
        X"1208812e",
        X"098106ff",
        X"9a38843d",
        X"0d04fe3d",
        X"0d805375",
        X"52745181",
        X"923f843d",
        X"0d04fe3d",
        X"0d815375",
        X"52745181",
        X"823f843d",
        X"0d04fb3d",
        X"0d777955",
        X"55805674",
        X"76258638",
        X"74305581",
        X"56738025",
        X"88387330",
        X"76813257",
        X"54805373",
        X"52745180",
        X"d63f83e0",
        X"80085475",
        X"802e8738",
        X"83e08008",
        X"30547383",
        X"e0800c87",
        X"3d0d04fa",
        X"3d0d787a",
        X"57558057",
        X"74772586",
        X"38743055",
        X"8157759f",
        X"2c548153",
        X"75743274",
        X"31527451",
        X"9a3f83e0",
        X"80085476",
        X"802e8738",
        X"83e08008",
        X"30547383",
        X"e0800c88",
        X"3d0d04fc",
        X"3d0d7678",
        X"53548153",
        X"80558739",
        X"71107310",
        X"54527372",
        X"26517280",
        X"2ea73870",
        X"802e8638",
        X"718025e8",
        X"3872802e",
        X"98387174",
        X"26893873",
        X"72317574",
        X"07565472",
        X"812a7281",
        X"2a5353e5",
        X"39735178",
        X"83387451",
        X"7083e080",
        X"0c863d0d",
        X"04fd3d0d",
        X"75775452",
        X"80547181",
        X"06ff1170",
        X"09750616",
        X"74812a76",
        X"10575556",
        X"515171ea",
        X"387383e0",
        X"800c853d",
        X"0d04fd3d",
        X"0d757771",
        X"ff1b5456",
        X"545270ff",
        X"2e923872",
        X"70810554",
        X"33727081",
        X"055434ff",
        X"1151eb39",
        X"7383e080",
        X"0c853d0d",
        X"04000000",
        X"00ffffff",
        X"ff00ffff",
        X"ffff00ff",
        X"ffffff00",
        X"809a9041",
        X"8e418f80",
        X"45454549",
        X"49498e8f",
        X"9092924f",
        X"994f5555",
        X"59999a9b",
        X"9c9d9e9f",
        X"41494f55",
        X"a5a5a6a7",
        X"a8a9aaab",
        X"ac21aeaf",
        X"b0b1b2b3",
        X"b4b5b6b7",
        X"b8b9babb",
        X"bcbdbebf",
        X"c0c1c2c3",
        X"c4c5c6c7",
        X"c8c9cacb",
        X"cccdcecf",
        X"d0d1d2d3",
        X"d4d5d6d7",
        X"d8d9dadb",
        X"dcdddedf",
        X"e0e1e2e3",
        X"e4e5e6e7",
        X"e8e9eaeb",
        X"ecedeeef",
        X"f0f1f2f3",
        X"f4f5f6f7",
        X"f8f9fafb",
        X"fcfdfeff",
        X"00000000",
        X"70704740",
        X"2c704268",
        X"2c020202",
        X"02020202",
        X"02020202",
        X"02020202",
        X"02020202",
        X"02020241",
        X"00060000",
        X"00002e8f",
        X"00002ed0",
        X"00002ef5",
        X"00002f07",
        X"00002f1b",
        X"2e2e0000",
        X"41545200",
        X"58464400",
        X"58455800",
        X"43686f6f",
        X"73652000",
        X"66696c65",
        X"00000000",
        X"4449523a",
        X"00000000",
        X"44495200",
        X"25732025",
        X"73000000",
        X"20000000",
        X"25303278",
        X"00000000",
        X"556e6b6e",
        X"6f776e20",
        X"74797065",
        X"206f6620",
        X"63617274",
        X"72696467",
        X"65210000",
        X"41353200",
        X"43415200",
        X"42494e00",
        X"31366b20",
        X"63617274",
        X"20747970",
        X"65000000",
        X"4c656674",
        X"20666f72",
        X"206f6e65",
        X"20636869",
        X"70000000",
        X"52696768",
        X"7420666f",
        X"72207477",
        X"6f206368",
        X"69700000",
        X"53650000",
        X"7474696e",
        X"67730000",
        X"54757262",
        X"6f3a2564",
        X"78000000",
        X"526f6d3a",
        X"25730000",
        X"4e4f4e45",
        X"00000000",
        X"43617274",
        X"3a257300",
        X"343a3300",
        X"31363a39",
        X"00000000",
        X"41737065",
        X"63742052",
        X"6174696f",
        X"3a202573",
        X"00000000",
        X"45786974",
        X"00000000",
        X"35323030",
        X"2e726f6d",
        X"00000000",
        X"524f4d00",
        X"4d454d00",
        X"00000000",
        X"00000000",
        X"01010008",
        X"02210010",
        X"080d0040",
        X"090a0040",
        X"0a090040",
        X"0b080040",
        X"0c300020",
        X"0d310040",
        X"0e320080",
        X"0f040010",
        X"110c0080",
        X"17330100",
        X"18340200",
        X"1a280010",
        X"1b290020",
        X"1c2a0040",
        X"1d2b0080",
        X"1e2c0100",
        X"1f2d0200",
        X"21380020",
        X"22390040",
        X"233a0080",
        X"243b0100",
        X"253c0200",
        X"28230010",
        X"29020080",
        X"2a030400",
        X"38240200",
        X"00000000",
        X"00000000",
        X"2f617461",
        X"72353230",
        X"302f726f",
        X"6d000000",
        X"2f617461",
        X"72353230",
        X"302f7573",
        X"65720000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000",
        X"00000000"

);

signal rdata:std_logic_vector(31 downto 0);
begin
        rdata<=ROM(conv_integer(address));

        process(clock)
        begin
                if(clock'event and clock='1')then
                	q<=rdata;
                end if;
        end process;
end syn;
